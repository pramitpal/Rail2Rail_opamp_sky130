magic
tech sky130A
magscale 1 2
timestamp 1678628286
<< nwell >>
rect 392 1992 1948 2008
rect 2472 1992 2782 1996
rect -446 1724 46 1726
rect 392 1724 2782 1992
rect -708 1688 2782 1724
rect -708 50 648 1688
rect 1720 449 2782 1688
rect 1720 448 2602 449
rect 2607 448 2782 449
rect 1720 398 2782 448
rect 1718 266 2782 398
rect 1718 116 2502 266
rect 1718 108 2484 116
rect 2488 108 2502 116
rect 1718 -12 2502 108
<< psubdiff >>
rect 1362 -1500 2090 -1480
rect 1362 -1506 1896 -1500
rect 1362 -1580 1396 -1506
rect 1548 -1574 1896 -1506
rect 2048 -1574 2090 -1500
rect 1548 -1580 2090 -1574
rect 1362 -1602 2090 -1580
<< nsubdiff >>
rect 706 1910 1486 1936
rect 706 1828 750 1910
rect 958 1908 1486 1910
rect 958 1828 1214 1908
rect 1442 1828 1486 1908
rect 706 1810 1486 1828
<< psubdiffcont >>
rect 1396 -1580 1548 -1506
rect 1896 -1574 2048 -1500
<< nsubdiffcont >>
rect 750 1828 958 1910
rect 1214 1828 1442 1908
<< poly >>
rect -288 1083 -202 1170
rect -288 1073 -87 1083
rect -288 1007 -169 1073
rect -103 1007 -87 1073
rect -288 997 -87 1007
rect 1956 796 2036 812
rect 1954 734 2036 796
rect 1950 724 2042 734
rect 1950 664 1966 724
rect 2026 710 2042 724
rect 2154 710 2234 810
rect 2026 664 2234 710
rect 1950 654 2234 664
rect 1956 630 2234 654
rect 2523 400 2589 407
rect 2648 400 2688 444
rect 2523 397 2688 400
rect 2523 363 2539 397
rect 2573 363 2688 397
rect 2523 360 2688 363
rect 2523 353 2589 360
rect 2484 258 2678 298
rect 2498 173 2538 258
rect 2638 206 2678 258
rect 2491 157 2545 173
rect -546 49 -436 124
rect -546 -22 -536 49
rect -446 -22 -436 49
rect -546 -38 -436 -22
rect -350 29 -240 104
rect -350 -42 -340 29
rect -250 -42 -240 29
rect -350 -58 -240 -42
rect 130 -26 248 62
rect 130 -32 299 -26
rect 398 -32 498 62
rect 848 54 908 122
rect 848 14 858 54
rect 898 14 908 54
rect 1204 22 1264 128
rect 2491 123 2501 157
rect 2535 123 2545 157
rect 2491 107 2545 123
rect 2296 61 2328 62
rect 848 -2 908 14
rect 1198 12 1270 22
rect 130 -42 498 -32
rect 1198 -28 1214 12
rect 1254 -28 1270 12
rect 1198 -38 1270 -28
rect 1906 9 1978 48
rect 2033 9 2103 15
rect 2296 9 2373 61
rect 1906 -1 2373 9
rect 130 -76 255 -42
rect 289 -76 498 -42
rect 1906 -51 2043 -1
rect 2093 -51 2373 -1
rect 1906 -61 2373 -51
rect 2033 -67 2103 -61
rect 130 -86 498 -76
rect 245 -92 299 -86
rect 368 -136 468 -129
rect 178 -139 468 -136
rect 178 -140 408 -139
rect 106 -206 408 -140
rect 106 -270 182 -206
rect 368 -213 408 -206
rect 452 -213 468 -139
rect 368 -216 468 -213
rect 368 -280 462 -216
rect 2060 -249 2263 -239
rect 2060 -278 2175 -249
rect 2056 -287 2175 -278
rect 2213 -287 2263 -249
rect 2056 -297 2263 -287
rect 2056 -354 2118 -297
rect 2060 -368 2118 -354
rect 2205 -365 2263 -297
rect 206 -1288 306 -1208
rect 364 -1288 464 -1204
rect 206 -1364 464 -1288
rect 1058 -1292 1122 -1288
rect 722 -1364 786 -1358
rect 1058 -1364 1130 -1292
rect 206 -1374 1130 -1364
rect 206 -1418 732 -1374
rect 776 -1388 1130 -1374
rect 776 -1418 1122 -1388
rect 206 -1424 1122 -1418
rect 428 -1428 1122 -1424
rect 722 -1434 786 -1428
<< polycont >>
rect -169 1007 -103 1073
rect 1966 664 2026 724
rect 2539 363 2573 397
rect -536 -22 -446 49
rect -340 -42 -250 29
rect 858 14 898 54
rect 2501 123 2535 157
rect 1214 -28 1254 12
rect 255 -76 289 -42
rect 2043 -51 2093 -1
rect 408 -213 452 -139
rect 2175 -287 2213 -249
rect 732 -1418 776 -1374
<< locali >>
rect 706 1910 1486 1934
rect 706 1828 750 1910
rect 958 1908 1486 1910
rect 958 1904 1214 1908
rect 958 1834 982 1904
rect 1198 1834 1214 1904
rect 958 1828 1214 1834
rect 1442 1828 1486 1908
rect 706 1808 1486 1828
rect -169 1073 -103 1089
rect -103 1013 -9 1067
rect -169 991 -103 1007
rect -552 -22 -536 49
rect -445 -22 -430 49
rect -356 -42 -340 29
rect -249 -42 -234 29
rect -63 -843 -9 1013
rect 1966 734 2026 740
rect 1676 724 2036 734
rect 1676 720 1966 724
rect 1744 664 1966 720
rect 2026 664 2036 724
rect 1744 654 2036 664
rect 1744 648 1772 654
rect 1966 648 2026 654
rect 2539 400 2573 413
rect 2539 347 2573 360
rect 2485 123 2498 157
rect 2538 123 2551 157
rect 842 14 848 54
rect 908 14 914 54
rect 1214 22 1254 28
rect 2033 -1 2103 9
rect 239 -76 245 -42
rect 299 -76 305 -42
rect 1214 -44 1254 -38
rect 2027 -51 2043 -1
rect 2093 -51 2109 -1
rect 408 -139 452 -123
rect 398 -208 408 -144
rect 452 -180 684 -144
rect 2033 -180 2103 -51
rect 452 -208 2103 -180
rect 408 -229 452 -213
rect 620 -209 2103 -208
rect 620 -238 2100 -209
rect 620 -242 684 -238
rect 2175 -239 2213 -233
rect 2175 -303 2213 -297
rect -63 -897 39 -843
rect 722 -1374 786 -1262
rect 716 -1418 732 -1374
rect 776 -1418 792 -1374
rect 722 -1428 786 -1418
rect 1362 -1496 2090 -1480
rect 1362 -1506 1628 -1496
rect 1362 -1580 1396 -1506
rect 1548 -1570 1628 -1506
rect 1780 -1500 2090 -1496
rect 1780 -1570 1896 -1500
rect 1548 -1574 1896 -1570
rect 2048 -1574 2090 -1500
rect 1548 -1580 2090 -1574
rect 1362 -1602 2090 -1580
<< viali >>
rect 982 1834 1198 1904
rect -536 49 -445 59
rect -536 -22 -446 49
rect -446 -22 -445 49
rect -340 29 -249 39
rect -536 -32 -445 -22
rect -340 -42 -250 29
rect -250 -42 -249 29
rect -340 -52 -249 -42
rect 1672 648 1744 720
rect 2536 397 2576 400
rect 2536 363 2539 397
rect 2539 363 2573 397
rect 2573 363 2576 397
rect 2536 360 2576 363
rect 2498 157 2538 160
rect 2498 123 2501 157
rect 2501 123 2535 157
rect 2535 123 2538 157
rect 2498 120 2538 123
rect 848 54 908 64
rect 848 14 858 54
rect 858 14 898 54
rect 898 14 908 54
rect 848 4 908 14
rect 1204 12 1264 22
rect 1204 -28 1214 12
rect 1214 -28 1254 12
rect 1254 -28 1264 12
rect 245 -42 299 -32
rect 1204 -38 1264 -28
rect 245 -76 255 -42
rect 255 -76 289 -42
rect 289 -76 299 -42
rect 245 -86 299 -76
rect 2165 -249 2223 -239
rect 2165 -287 2175 -249
rect 2175 -287 2213 -249
rect 2213 -287 2223 -249
rect 2165 -297 2223 -287
rect 39 -897 93 -843
rect 1628 -1570 1780 -1496
<< metal1 >>
rect 596 1904 1532 1972
rect -146 1784 -102 1904
rect 596 1834 982 1904
rect 1198 1834 1532 1904
rect 596 1784 1532 1834
rect -146 1783 2146 1784
rect -146 1740 2640 1783
rect -146 1566 -102 1740
rect 300 1620 344 1740
rect 2097 1730 2640 1740
rect 2100 1600 2146 1730
rect -406 894 -362 1232
rect 762 851 1877 880
rect 762 809 1883 851
rect 774 526 820 809
rect 1660 720 1756 726
rect 1290 674 1340 677
rect 1464 674 1470 685
rect 1290 630 1470 674
rect 1290 528 1340 630
rect 1464 620 1470 630
rect 1535 620 1541 685
rect 1660 648 1672 720
rect 1744 648 1756 720
rect 1660 642 1756 648
rect 690 408 742 414
rect 565 357 690 407
rect 690 350 742 356
rect -666 -503 -622 184
rect -548 59 -433 65
rect -548 53 -536 59
rect -445 53 -433 59
rect -548 -38 -542 53
rect -439 -38 -433 53
rect -352 39 -334 45
rect -542 -44 -439 -38
rect -352 -52 -340 39
rect -352 -58 -334 -52
rect -243 -58 -237 45
rect -666 -548 -282 -503
rect -140 -532 -96 148
rect 44 -82 88 102
rect 36 -83 88 -82
rect 233 -32 311 -26
rect 233 -83 245 -32
rect 36 -86 245 -83
rect 299 -86 311 -32
rect 36 -92 311 -86
rect 36 -132 299 -92
rect 36 -148 83 -132
rect 34 -298 83 -148
rect 558 -166 602 86
rect 836 64 920 70
rect 836 4 848 64
rect 908 4 920 64
rect 836 -2 920 4
rect 314 -210 602 -166
rect 314 -316 358 -210
rect 848 -346 908 -2
rect 1031 -109 1077 247
rect 1198 28 1270 34
rect 1192 -44 1198 28
rect 1258 22 1270 28
rect 1264 -38 1270 22
rect 1258 -44 1270 -38
rect 1198 -50 1270 -44
rect 578 -406 584 -346
rect 644 -406 838 -346
rect 898 -406 908 -346
rect 960 -155 1077 -109
rect 960 -522 1006 -155
rect -663 -549 -282 -548
rect -331 -721 -285 -549
rect -150 -584 -144 -532
rect -92 -584 -86 -532
rect 566 -584 572 -532
rect 624 -584 630 -532
rect 196 -705 238 -632
rect 155 -721 238 -705
rect -331 -747 238 -721
rect 474 -704 516 -652
rect 576 -704 620 -584
rect -331 -767 197 -747
rect 151 -805 197 -767
rect 474 -748 620 -704
rect 474 -798 516 -748
rect 27 -843 105 -837
rect 27 -897 39 -843
rect 93 -897 105 -843
rect 155 -847 197 -805
rect 27 -903 105 -897
rect 1672 -869 1744 642
rect 1837 595 1883 809
rect 2253 685 2318 691
rect 2253 597 2318 620
rect 2365 597 2411 847
rect 1837 549 2032 595
rect 1986 450 2032 549
rect 2244 551 2411 597
rect 2244 544 2318 551
rect 2244 462 2290 544
rect 2530 406 2582 412
rect 2524 354 2530 406
rect 2582 354 2588 406
rect 2530 348 2582 354
rect 2705 320 2751 523
rect 2705 319 2788 320
rect 2705 315 2772 319
rect 2686 269 2772 315
rect 2486 160 2550 166
rect 1819 -98 1865 127
rect 2486 120 2498 160
rect 2538 120 2550 160
rect 2686 148 2732 269
rect 2766 266 2772 269
rect 2825 266 2862 319
rect 2486 116 2550 120
rect 2488 114 2550 116
rect 2413 60 2459 87
rect 2498 60 2538 114
rect 2413 20 2538 60
rect 1819 -144 2004 -98
rect 1958 -239 2004 -144
rect 2413 -167 2459 20
rect 2298 -213 2459 -167
rect 2159 -239 2229 -227
rect 1958 -297 2165 -239
rect 2223 -297 2229 -239
rect 1958 -303 2031 -297
rect 1985 -419 2031 -303
rect 2159 -309 2229 -297
rect 2298 -384 2344 -213
rect 2140 -869 2186 -756
rect 39 -1110 93 -903
rect 1672 -915 2625 -869
rect 39 -1167 101 -1110
rect 55 -1439 101 -1167
rect 312 -1439 358 -1194
rect 55 -1440 358 -1439
rect 1218 -1440 1264 -1262
rect 1672 -1440 1744 -915
rect 55 -1442 1744 -1440
rect 55 -1485 2132 -1442
rect 312 -1486 2132 -1485
rect 1326 -1496 2132 -1486
rect 1326 -1570 1628 -1496
rect 1780 -1570 2132 -1496
rect 1326 -1634 2132 -1570
<< via1 >>
rect 1470 620 1535 685
rect 690 356 742 408
rect -542 -32 -536 53
rect -536 -32 -445 53
rect -445 -32 -439 53
rect -542 -38 -439 -32
rect -334 39 -243 45
rect -334 -52 -249 39
rect -249 -52 -243 39
rect -334 -58 -243 -52
rect 1198 22 1258 28
rect 1198 -38 1204 22
rect 1204 -38 1258 22
rect 1198 -44 1258 -38
rect 584 -406 644 -346
rect 838 -406 898 -346
rect -144 -584 -92 -532
rect 572 -584 624 -532
rect 2253 620 2318 685
rect 2530 400 2582 406
rect 2530 360 2536 400
rect 2536 360 2576 400
rect 2576 360 2582 400
rect 2530 354 2582 360
rect 2772 266 2825 319
<< metal2 >>
rect 1470 685 1535 691
rect 1535 620 2253 685
rect 2318 620 2324 685
rect 1470 614 1535 620
rect 684 356 690 408
rect 742 407 748 408
rect 742 405 2482 407
rect 2530 406 2582 412
rect 742 357 2530 405
rect 742 356 748 357
rect 2482 355 2530 357
rect 2530 348 2582 354
rect 2772 319 2825 325
rect 1480 266 2772 319
rect -548 -38 -542 53
rect -439 -38 -433 53
rect -334 45 -243 51
rect -535 -346 -444 -38
rect 1198 28 1258 34
rect -243 22 912 25
rect -243 -37 1198 22
rect 872 -38 1198 -37
rect 1198 -50 1258 -44
rect -334 -64 -243 -58
rect 584 -346 644 -340
rect -535 -406 584 -346
rect -535 -407 -444 -406
rect 584 -412 644 -406
rect 838 -346 898 -340
rect 1480 -346 1533 266
rect 2772 260 2825 266
rect 898 -406 1533 -346
rect 838 -412 898 -406
rect -144 -532 -92 -526
rect 572 -532 624 -526
rect -92 -580 572 -536
rect -144 -590 -92 -584
rect 572 -590 624 -584
use sky130_fd_pr__nfet_01v8_42C9PJ  sky130_fd_pr__nfet_01v8_42C9PJ_0
timestamp 1678605198
transform 1 0 2163 0 1 -568
box -187 -226 187 226
use sky130_fd_pr__nfet_01v8_42C9PJ  sky130_fd_pr__nfet_01v8_42C9PJ_1
timestamp 1678605198
transform 1 0 335 0 1 -998
box -187 -226 187 226
use sky130_fd_pr__nfet_01v8_C5U7X2  sky130_fd_pr__nfet_01v8_C5U7X2_0
timestamp 1678605198
transform 1 0 2658 0 1 -610
box -78 -826 78 826
use sky130_fd_pr__nfet_01v8_SAC9P4  sky130_fd_pr__nfet_01v8_SAC9P4_0
timestamp 1678605198
transform 1 0 414 0 1 -484
box -108 -226 108 226
use sky130_fd_pr__nfet_01v8_SAC9P4  sky130_fd_pr__nfet_01v8_SAC9P4_1
timestamp 1678605198
transform 1 0 136 0 1 -474
box -108 -226 108 226
use sky130_fd_pr__nfet_01v8_SLJEK5  sky130_fd_pr__nfet_01v8_SLJEK5_0
timestamp 1678603392
transform 1 0 1112 0 1 -888
box -158 -426 158 426
use sky130_fd_pr__nfet_01v8_VYPHSS  sky130_fd_pr__nfet_01v8_VYPHSS_0
timestamp 1678603392
transform 1 0 1055 0 1 336
box -287 -226 287 226
use sky130_fd_pr__pfet_01v8_7Q88LS  sky130_fd_pr__pfet_01v8_7Q88LS_0
timestamp 1678602466
transform 1 0 -383 0 1 516
box -323 -462 323 462
use sky130_fd_pr__pfet_01v8_7Q88LS  sky130_fd_pr__pfet_01v8_7Q88LS_1
timestamp 1678602466
transform 1 0 2123 0 1 1212
box -323 -462 323 462
use sky130_fd_pr__pfet_01v8_9Q4LM2  sky130_fd_pr__pfet_01v8_9Q4LM2_0
timestamp 1678601982
transform 1 0 -252 0 1 1382
box -194 -262 194 262
use sky130_fd_pr__pfet_01v8_EE9SH3  sky130_fd_pr__pfet_01v8_EE9SH3_0
timestamp 1678605198
transform 1 0 2668 0 1 1452
box -114 -1062 114 1062
use sky130_fd_pr__pfet_01v8_SK88LG  sky130_fd_pr__pfet_01v8_SK88LG_0
timestamp 1678601982
transform 1 0 323 0 1 862
box -323 -862 323 862
use sky130_fd_pr__pfet_01v8_W7GQZ7  sky130_fd_pr__pfet_01v8_W7GQZ7_0
timestamp 1678605484
transform 1 0 2346 0 1 264
box -144 -262 144 262
use sky130_fd_pr__pfet_01v8_W7GQZ7  sky130_fd_pr__pfet_01v8_W7GQZ7_1
timestamp 1678605484
transform 1 0 1928 0 1 260
box -144 -262 144 262
<< labels >>
flabel metal1 s -124 1864 -124 1864 0 FreeSans 800 0 0 0 VDD
port 1 nsew
flabel metal1 s 318 -1458 318 -1458 0 FreeSans 800 0 0 0 GND
port 3 nsew
flabel locali s 760 -1294 760 -1294 0 FreeSans 800 0 0 0 VB2
port 4 nsew
flabel metal2 s 1140 -6 1140 -6 0 FreeSans 800 0 0 0 PLUS
port 5 nsew
flabel metal1 s 2836 288 2836 288 0 FreeSans 800 0 0 0 OUT3
port 6 nsew
flabel locali s 674 -208 674 -208 1 FreeSans 1600 0 0 0 VB1
port 7 n
<< end >>
