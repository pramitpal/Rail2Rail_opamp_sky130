magic
tech sky130A
magscale 1 2
timestamp 1681052864
<< nwell >>
rect 677 3755 3685 3957
rect 697 2969 3685 3755
rect 1323 2691 3685 2969
rect 1323 2141 1832 2691
rect 1414 228 2112 1825
rect 2837 1707 3683 2691
rect 1423 226 2110 228
<< psubdiff >>
rect 27 123 1213 131
rect 27 30 87 123
rect 180 30 276 123
rect 369 30 450 123
rect 543 30 633 123
rect 726 30 820 123
rect 913 30 1023 123
rect 1116 30 1213 123
rect 27 22 1213 30
<< nsubdiff >>
rect 1202 3869 1886 3877
rect 1202 3756 1243 3869
rect 1333 3756 1404 3869
rect 1517 3756 1673 3869
rect 1786 3868 1886 3869
rect 1786 3860 2734 3868
rect 1786 3768 1967 3860
rect 2059 3768 2156 3860
rect 2248 3768 2350 3860
rect 2442 3768 2555 3860
rect 2647 3768 2734 3860
rect 1786 3760 2734 3768
rect 1786 3756 1886 3760
rect 1202 3748 1886 3756
<< psubdiffcont >>
rect 87 30 180 123
rect 276 30 369 123
rect 450 30 543 123
rect 633 30 726 123
rect 820 30 913 123
rect 1023 30 1116 123
<< nsubdiffcont >>
rect 1243 3756 1333 3869
rect 1404 3756 1517 3869
rect 1673 3756 1786 3869
rect 1967 3768 2059 3860
rect 2156 3768 2248 3860
rect 2350 3768 2442 3860
rect 2555 3768 2647 3860
<< poly >>
rect 1230 3121 1284 3134
rect 1480 3121 1520 3147
rect 1230 3118 1520 3121
rect 1230 3084 1240 3118
rect 1274 3084 1520 3118
rect 1230 3081 1520 3084
rect 1230 3068 1284 3081
rect 716 2935 770 2950
rect 854 2935 891 3030
rect 1012 2944 1049 3035
rect 986 2935 1052 2944
rect 716 2934 1052 2935
rect 716 2900 726 2934
rect 760 2900 1002 2934
rect 1036 2900 1052 2934
rect 716 2898 1052 2900
rect 716 2884 770 2898
rect 986 2890 1052 2898
rect 940 2818 1006 2828
rect 940 2784 956 2818
rect 990 2784 1006 2818
rect 940 2774 1006 2784
rect 958 2732 988 2774
rect 958 2722 992 2732
rect 958 2702 988 2722
rect 2258 2647 2304 2798
rect 2248 2643 2314 2647
rect 2421 2643 2467 2788
rect 2248 2637 2467 2643
rect 2248 2603 2264 2637
rect 2298 2603 2467 2637
rect 2248 2597 2467 2603
rect 2248 2593 2314 2597
rect 1478 2063 1518 2214
rect 1638 2064 1675 2213
rect 1471 2047 1525 2063
rect 1471 2013 1481 2047
rect 1515 2013 1525 2047
rect 1471 1997 1525 2013
rect 1630 2048 1684 2064
rect 1630 2014 1640 2048
rect 1674 2014 1684 2048
rect 1630 1998 1684 2014
rect 2203 2044 2246 2124
rect 2483 2044 2526 2125
rect 2203 2001 2693 2044
rect 2650 1895 2693 2001
rect 2645 1879 2699 1895
rect 1014 1845 1068 1861
rect 1014 1811 1024 1845
rect 1058 1811 1068 1845
rect 1014 1795 1068 1811
rect 1177 1841 1231 1857
rect 1177 1807 1187 1841
rect 1221 1807 1231 1841
rect 1020 1713 1062 1795
rect 1177 1791 1231 1807
rect 2337 1842 2391 1858
rect 2337 1808 2347 1842
rect 2381 1808 2391 1842
rect 2645 1845 2655 1879
rect 2689 1845 2699 1879
rect 2645 1829 2699 1845
rect 2337 1798 2391 1808
rect 1184 1715 1223 1791
rect 2274 1758 2457 1798
rect 2274 1682 2314 1758
rect 2417 1683 2457 1758
rect 1662 831 1712 953
rect 1814 831 1864 937
rect 1379 781 1864 831
rect 1379 720 1429 781
rect 2280 770 2346 778
rect 2280 768 2626 770
rect 2280 734 2296 768
rect 2330 734 2626 768
rect 2280 731 2626 734
rect 2280 724 2346 731
rect 1371 710 1437 720
rect 1371 676 1387 710
rect 1421 676 1437 710
rect 1371 666 1437 676
rect 2423 585 2462 731
rect 2587 590 2626 731
rect 1033 259 1073 383
rect 1026 243 1080 259
rect 1026 209 1036 243
rect 1070 209 1080 243
rect 1026 193 1080 209
rect 1351 208 1417 218
rect 1584 208 1618 298
rect 1929 208 1963 297
rect 2113 208 2179 218
rect 1351 174 1367 208
rect 1401 174 2129 208
rect 2163 174 2179 208
rect 1351 164 1417 174
rect 2113 164 2179 174
<< polycont >>
rect 1240 3084 1274 3118
rect 726 2900 760 2934
rect 1002 2900 1036 2934
rect 956 2784 990 2818
rect 2264 2603 2298 2637
rect 1481 2013 1515 2047
rect 1640 2014 1674 2048
rect 1024 1811 1058 1845
rect 1187 1807 1221 1841
rect 2347 1808 2381 1842
rect 2655 1845 2689 1879
rect 2296 734 2330 768
rect 1387 676 1421 710
rect 1036 209 1070 243
rect 1367 174 1401 208
rect 2129 174 2163 208
<< locali >>
rect 1862 3900 2788 3933
rect 1172 3869 2788 3900
rect 1172 3756 1243 3869
rect 1333 3866 1404 3869
rect 1517 3863 1673 3869
rect 1333 3756 1404 3773
rect 1517 3766 1544 3863
rect 1644 3766 1673 3863
rect 1517 3756 1673 3766
rect 1786 3862 2788 3869
rect 1786 3860 2530 3862
rect 1786 3858 1967 3860
rect 2059 3859 2156 3860
rect 1786 3765 1799 3858
rect 1876 3768 1967 3858
rect 2248 3857 2350 3860
rect 2248 3768 2271 3857
rect 2442 3770 2530 3860
rect 2651 3770 2788 3862
rect 2967 3875 3596 3923
rect 2919 3783 2967 3875
rect 3234 3778 3282 3875
rect 3548 3846 3596 3875
rect 3548 3823 3598 3846
rect 3550 3778 3598 3823
rect 2442 3768 2555 3770
rect 2647 3768 2788 3770
rect 1876 3767 2036 3768
rect 2157 3767 2271 3768
rect 1876 3765 2271 3767
rect 2392 3765 2788 3768
rect 1786 3756 2788 3765
rect 1172 3718 2788 3756
rect 1862 3717 2788 3718
rect 775 3022 812 3088
rect 725 2985 812 3022
rect 725 2950 762 2985
rect 660 2934 770 2950
rect 1002 2936 1036 2950
rect 660 2900 726 2934
rect 760 2900 776 2934
rect 660 2867 770 2900
rect 1002 2884 1036 2899
rect 660 1359 724 2867
rect 956 2818 990 2834
rect 1095 2818 1129 3129
rect 1224 3084 1237 3118
rect 1277 3084 1290 3118
rect 990 2784 1129 2818
rect 956 2768 990 2784
rect 1038 2719 1072 2784
rect 1037 2704 1072 2719
rect 1037 2703 1071 2704
rect 1040 2691 1069 2703
rect 2171 2643 2217 2879
rect 2264 2643 2298 2653
rect 2171 2637 2304 2643
rect 2171 2603 2264 2637
rect 2298 2603 2304 2637
rect 2658 2606 2783 2651
rect 2670 2604 2783 2606
rect 2171 2597 2304 2603
rect 2264 2587 2298 2597
rect 1030 2146 1067 2509
rect 2736 2369 2783 2604
rect 1725 2258 2048 2301
rect 1030 2106 1918 2146
rect 1030 2076 1067 2106
rect 0 1293 110 1354
rect 542 1276 724 1359
rect 765 2039 1067 2076
rect 1478 2047 1518 2050
rect 1639 2048 1676 2050
rect 163 990 567 993
rect 163 956 530 990
rect 564 956 567 990
rect 163 954 567 956
rect 619 713 669 1276
rect 619 675 624 713
rect 664 675 669 713
rect 619 669 669 675
rect 185 306 682 340
rect 765 244 802 2039
rect 1465 2013 1481 2047
rect 1515 2013 1531 2047
rect 1624 2014 1640 2048
rect 1674 2014 1690 2048
rect 1478 1958 1518 2013
rect 1020 1920 1415 1958
rect 1453 1920 1518 1958
rect 1020 1918 1518 1920
rect 1020 1882 1060 1918
rect 1639 1884 1676 2014
rect 1020 1845 1062 1882
rect 1185 1845 1676 1884
rect 1878 1903 1918 2106
rect 2005 2029 2048 2258
rect 2005 2024 2560 2029
rect 2005 1990 2521 2024
rect 2555 1990 2560 2024
rect 2005 1986 2560 1990
rect 2834 1913 2883 1919
rect 2344 1903 2384 1904
rect 1878 1863 2384 1903
rect 2651 1879 2694 1884
rect 1008 1811 1024 1845
rect 1058 1811 1074 1845
rect 1185 1841 1237 1845
rect 1020 1807 1062 1811
rect 1171 1807 1187 1841
rect 1221 1807 1237 1841
rect 1185 1805 1224 1807
rect 1366 1446 1405 1845
rect 2331 1842 2384 1863
rect 2639 1845 2655 1879
rect 2689 1845 2705 1879
rect 2834 1876 2840 1913
rect 2877 1876 2883 1913
rect 2331 1808 2347 1842
rect 2381 1808 2397 1842
rect 2344 1805 2384 1808
rect 2651 1246 2694 1845
rect 2834 1676 2883 1876
rect 2834 1665 3613 1676
rect 2730 1662 3613 1665
rect 2730 1628 2733 1662
rect 2767 1628 3613 1662
rect 2730 1627 3613 1628
rect 2730 1625 2873 1627
rect 2114 1203 2694 1246
rect 1312 853 1361 1145
rect 1312 846 1878 853
rect 1312 809 1835 846
rect 1872 809 1878 846
rect 1312 804 1878 809
rect 1387 718 1421 726
rect 1387 660 1421 668
rect 876 244 1073 246
rect 765 243 1073 244
rect 765 209 1036 243
rect 1070 209 1086 243
rect 2114 226 2157 1203
rect 2208 771 2260 774
rect 2296 771 2330 784
rect 2208 768 2333 771
rect 2208 734 2296 768
rect 2330 734 2333 768
rect 2208 732 2333 734
rect 2208 594 2260 732
rect 2296 718 2330 732
rect 2807 713 2850 1520
rect 2373 708 2850 713
rect 2373 674 2377 708
rect 2411 674 2850 708
rect 2373 670 2850 674
rect 2208 542 2389 594
rect 2665 535 2708 670
rect 765 207 1073 209
rect 1367 208 1401 224
rect 876 206 1073 207
rect 1331 174 1367 208
rect 1367 158 1401 174
rect 2114 208 2186 226
rect 2114 174 2129 208
rect 2163 174 2186 208
rect 2114 164 2186 174
rect 2117 157 2186 164
rect 2805 177 2845 310
rect 3084 177 3124 322
rect 3402 177 3442 313
rect 0 135 1251 157
rect 2805 137 3442 177
rect 0 131 722 135
rect 0 26 37 131
rect 141 129 543 131
rect 141 123 205 129
rect 309 123 374 129
rect 478 123 543 129
rect 647 123 722 131
rect 826 123 909 135
rect 1013 133 1251 135
rect 1013 123 1110 133
rect 180 30 205 123
rect 369 30 374 123
rect 1013 30 1023 123
rect 141 26 205 30
rect 0 24 205 26
rect 309 24 374 30
rect 478 26 543 30
rect 647 28 1110 30
rect 1214 28 1251 133
rect 647 26 1251 28
rect 478 24 1251 26
rect 0 0 1251 24
<< viali >>
rect 1332 3773 1333 3866
rect 1333 3773 1404 3866
rect 1404 3773 1409 3866
rect 1544 3766 1644 3863
rect 2530 3860 2651 3862
rect 1799 3765 1876 3858
rect 2036 3768 2059 3859
rect 2059 3768 2156 3859
rect 2156 3768 2157 3859
rect 2271 3768 2350 3857
rect 2350 3768 2392 3857
rect 2530 3770 2555 3860
rect 2555 3770 2647 3860
rect 2647 3770 2651 3860
rect 2919 3875 2967 3923
rect 2036 3767 2157 3768
rect 2271 3765 2392 3768
rect 1001 2934 1038 2936
rect 1001 2900 1002 2934
rect 1002 2900 1036 2934
rect 1036 2900 1038 2934
rect 1001 2899 1038 2900
rect 1237 3118 1277 3121
rect 1237 3084 1240 3118
rect 1240 3084 1274 3118
rect 1274 3084 1277 3118
rect 1237 3081 1277 3084
rect 2613 2606 2658 2651
rect 2736 2322 2783 2369
rect 110 1293 171 1354
rect 530 956 564 990
rect 624 675 664 713
rect 682 303 716 343
rect 1415 1920 1453 1958
rect 2521 1990 2555 2024
rect 2840 1876 2877 1913
rect 1366 1407 1405 1446
rect 2733 1628 2767 1662
rect 3613 1627 3662 1676
rect 2807 1520 2850 1563
rect 1312 1145 1361 1194
rect 1835 809 1872 846
rect 1379 710 1429 718
rect 1379 676 1387 710
rect 1387 676 1421 710
rect 1421 676 1429 710
rect 1379 668 1429 676
rect 2377 674 2411 708
rect 2805 310 2845 350
rect 1297 174 1331 208
rect 37 123 141 131
rect 205 123 309 129
rect 374 123 478 129
rect 543 123 647 131
rect 722 123 826 135
rect 909 123 1013 135
rect 1110 123 1214 133
rect 37 30 87 123
rect 87 30 141 123
rect 205 30 276 123
rect 276 30 309 123
rect 374 30 450 123
rect 450 30 478 123
rect 543 30 633 123
rect 633 30 647 123
rect 722 30 726 123
rect 726 30 820 123
rect 820 30 826 123
rect 909 30 913 123
rect 913 30 1013 123
rect 1110 30 1116 123
rect 1116 30 1214 123
rect 37 26 141 30
rect 205 24 309 30
rect 374 24 478 30
rect 543 26 647 30
rect 1110 28 1214 30
<< metal1 >>
rect 1862 3932 2788 3933
rect 931 3923 2788 3932
rect 2913 3923 2973 3935
rect 931 3885 2919 3923
rect 931 3811 978 3885
rect 1166 3875 2919 3885
rect 2967 3875 2973 3923
rect 1166 3866 2788 3875
rect 1166 3773 1332 3866
rect 1409 3863 2788 3866
rect 2913 3863 2973 3875
rect 3068 3872 3074 3924
rect 3126 3875 3445 3924
rect 3126 3872 3132 3875
rect 1409 3773 1544 3863
rect 1166 3766 1544 3773
rect 1644 3862 2788 3863
rect 1644 3859 2530 3862
rect 1644 3858 2036 3859
rect 1644 3766 1799 3858
rect 1166 3765 1799 3766
rect 1876 3767 2036 3858
rect 2157 3857 2530 3859
rect 2157 3767 2271 3857
rect 1876 3765 2271 3767
rect 2392 3770 2530 3857
rect 2651 3770 2788 3862
rect 3075 3796 3124 3872
rect 3392 3800 3441 3875
rect 2392 3765 2788 3770
rect 1166 3718 2788 3765
rect 1390 3522 1443 3718
rect 1862 3717 2788 3718
rect 1225 3121 1289 3127
rect 1225 3081 1237 3121
rect 1277 3081 1289 3121
rect 1225 3075 1289 3081
rect 995 2937 1044 2948
rect 1237 2937 1277 3075
rect 1557 2989 1605 3165
rect 995 2936 1277 2937
rect 995 2899 1001 2936
rect 1038 2900 1277 2936
rect 1038 2899 1044 2900
rect 995 2887 1044 2899
rect 1866 2399 1910 3717
rect 2331 3541 2378 3717
rect 2826 3620 2832 3672
rect 2884 3620 2890 3672
rect 2174 2676 2219 2834
rect 2174 2631 2322 2676
rect 2277 2483 2322 2631
rect 2505 2652 2550 2831
rect 2607 2652 2664 2663
rect 2505 2651 2664 2652
rect 2505 2627 2613 2651
rect 2392 2607 2613 2627
rect 2392 2582 2550 2607
rect 2607 2606 2613 2607
rect 2658 2606 2664 2651
rect 2607 2594 2664 2606
rect 2392 2484 2437 2582
rect 861 2171 922 2396
rect 1856 2347 1862 2399
rect 1914 2347 1920 2399
rect 2724 2369 2795 2375
rect 2724 2322 2736 2369
rect 2783 2322 2795 2369
rect 2724 2316 2795 2322
rect 745 2117 922 2171
rect 745 2110 921 2117
rect 745 1628 806 2110
rect 1383 2084 1426 2257
rect 1383 2078 1897 2084
rect 1383 2041 2048 2078
rect 1789 2040 2048 2041
rect 2118 2040 2161 2162
rect 1789 2035 2235 2040
rect 2005 1997 2235 2035
rect 2557 2030 2600 2154
rect 1784 1983 1836 1989
rect 1403 1958 1465 1964
rect 1403 1920 1415 1958
rect 1453 1920 1465 1958
rect 1403 1914 1465 1920
rect 1740 1931 1784 1936
rect 1740 1925 1836 1931
rect 412 1567 806 1628
rect 1409 1624 1459 1914
rect 1740 1892 1832 1925
rect 1740 1712 1784 1892
rect 2192 1645 2235 1997
rect 2509 2024 2600 2030
rect 2509 1990 2521 2024
rect 2555 1990 2600 2024
rect 2509 1985 2600 1990
rect 2509 1984 2567 1985
rect 2512 1654 2555 1984
rect 2736 1773 2783 2316
rect 2834 1913 2883 3620
rect 2834 1876 2840 1913
rect 2877 1876 2883 1913
rect 2834 1864 2883 1876
rect 2736 1726 3542 1773
rect 2951 1718 3542 1726
rect 3574 1676 3699 1703
rect 2721 1662 2779 1668
rect 2582 1624 2634 1630
rect 1402 1572 1408 1624
rect 1460 1572 1466 1624
rect 2721 1628 2733 1662
rect 2767 1628 2779 1662
rect 2721 1623 2779 1628
rect 2634 1622 2779 1623
rect 3574 1627 3613 1676
rect 3662 1627 3699 1676
rect 2634 1573 2770 1622
rect 3574 1596 3699 1627
rect 104 1355 177 1366
rect 412 1355 473 1567
rect 2582 1566 2634 1572
rect 835 1454 887 1460
rect 670 1409 835 1448
rect 104 1354 479 1355
rect 104 1293 110 1354
rect 171 1339 479 1354
rect 171 1294 481 1339
rect 171 1293 177 1294
rect 104 1281 177 1293
rect 435 157 481 1294
rect 518 992 576 996
rect 670 992 709 1409
rect 1360 1453 1411 1458
rect 835 1396 887 1402
rect 1354 1401 1360 1453
rect 1412 1401 1418 1453
rect 1360 1395 1411 1401
rect 937 1282 986 1376
rect 842 1233 986 1282
rect 842 1193 891 1233
rect 834 1141 840 1193
rect 892 1141 898 1193
rect 1106 1158 1154 1356
rect 2730 1340 2770 1573
rect 2801 1563 2856 1575
rect 2970 1563 3561 1565
rect 2801 1520 2807 1563
rect 2850 1520 3561 1563
rect 2801 1508 2856 1520
rect 2970 1510 3561 1520
rect 1259 1277 1305 1332
rect 1259 1231 1364 1277
rect 1312 1200 1361 1231
rect 1300 1194 1373 1200
rect 1300 1145 1312 1194
rect 1361 1145 1373 1194
rect 1300 1139 1373 1145
rect 2343 1063 2393 1307
rect 2730 1300 2845 1340
rect 2343 1013 2551 1063
rect 2343 1009 2393 1013
rect 518 990 709 992
rect 518 956 530 990
rect 564 956 709 990
rect 518 953 709 956
rect 518 950 576 953
rect 1285 917 1337 923
rect 1576 915 1625 986
rect 1337 866 1625 915
rect 1285 859 1337 865
rect 1576 846 1625 866
rect 1892 852 1941 965
rect 1823 846 1941 852
rect 1576 797 1702 846
rect 1823 809 1835 846
rect 1872 809 1941 846
rect 1823 803 1941 809
rect 618 719 670 725
rect 1373 724 1435 730
rect 612 667 618 719
rect 670 667 676 719
rect 618 663 670 667
rect 1367 662 1373 724
rect 1425 718 1435 724
rect 1429 668 1435 718
rect 1653 676 1702 797
rect 1829 684 1878 803
rect 2365 712 2423 714
rect 2216 708 2423 712
rect 1425 662 1435 668
rect 1373 656 1435 662
rect 2216 674 2377 708
rect 2411 674 2423 708
rect 2216 669 2423 674
rect 676 349 728 355
rect 670 297 676 349
rect 676 291 728 297
rect 947 157 993 386
rect 1291 217 1337 220
rect 1282 165 1288 217
rect 1340 165 1346 217
rect 1291 162 1337 165
rect 0 135 1251 157
rect 0 131 722 135
rect 0 26 37 131
rect 141 129 543 131
rect 141 26 205 129
rect 0 24 205 26
rect 309 24 374 129
rect 478 26 543 129
rect 647 30 722 131
rect 826 30 909 135
rect 1013 133 1251 135
rect 1013 30 1110 133
rect 647 28 1110 30
rect 1214 129 1251 133
rect 1494 150 1532 355
rect 1996 290 2072 338
rect 2216 290 2259 669
rect 2365 668 2423 669
rect 2501 538 2551 1013
rect 2805 356 2845 1300
rect 2793 350 2857 356
rect 2793 310 2805 350
rect 2845 310 2857 350
rect 2793 304 2857 310
rect 1996 247 2259 290
rect 2925 286 2972 287
rect 2348 150 2386 253
rect 1214 75 1260 129
rect 1494 112 2386 150
rect 2507 75 2553 256
rect 2925 255 2978 286
rect 2932 201 2978 255
rect 3246 201 3292 320
rect 3561 201 3607 335
rect 2932 155 3607 201
rect 2932 75 2978 155
rect 1214 29 2978 75
rect 1214 28 1260 29
rect 647 26 1260 28
rect 478 24 1260 26
rect 0 0 1260 24
<< via1 >>
rect 3074 3872 3126 3924
rect 2832 3620 2884 3672
rect 1862 2347 1914 2399
rect 1784 1931 1836 1983
rect 1408 1572 1460 1624
rect 2582 1572 2634 1624
rect 835 1402 887 1454
rect 1360 1446 1412 1453
rect 1360 1407 1366 1446
rect 1366 1407 1405 1446
rect 1405 1407 1412 1446
rect 1360 1401 1412 1407
rect 840 1141 892 1193
rect 1285 865 1337 917
rect 618 713 670 719
rect 618 675 624 713
rect 624 675 664 713
rect 664 675 670 713
rect 618 667 670 675
rect 1373 718 1425 724
rect 1373 668 1379 718
rect 1379 668 1425 718
rect 1373 662 1425 668
rect 676 343 728 349
rect 676 303 682 343
rect 682 303 716 343
rect 716 303 728 343
rect 676 297 728 303
rect 1288 208 1340 217
rect 1288 174 1297 208
rect 1297 174 1331 208
rect 1331 174 1340 208
rect 1288 165 1340 174
<< metal2 >>
rect 3074 3924 3126 3930
rect 2833 3874 3074 3923
rect 2833 3678 2882 3874
rect 3074 3866 3126 3872
rect 2832 3672 2884 3678
rect 2832 3614 2884 3620
rect 1862 2399 1914 2405
rect 1788 2351 1862 2395
rect 1788 1983 1832 2351
rect 1862 2341 1914 2347
rect 1778 1931 1784 1983
rect 1836 1931 1842 1983
rect 1408 1624 1460 1630
rect 1405 1573 1408 1623
rect 2576 1623 2582 1624
rect 1460 1573 2582 1623
rect 2576 1572 2582 1573
rect 2634 1572 2640 1624
rect 1408 1566 1460 1572
rect 829 1402 835 1454
rect 887 1447 893 1454
rect 1360 1453 1412 1459
rect 887 1408 1360 1447
rect 887 1402 893 1408
rect 1360 1395 1412 1401
rect 840 1193 892 1199
rect 892 1189 1328 1191
rect 892 1142 1336 1189
rect 840 1135 892 1141
rect 1287 917 1336 1142
rect 1279 865 1285 917
rect 1337 865 1343 917
rect 618 719 670 725
rect 1373 724 1425 730
rect 670 668 1373 718
rect 618 661 670 667
rect 1373 656 1425 662
rect 670 297 676 349
rect 728 297 734 349
rect 685 208 719 297
rect 1288 217 1340 223
rect 685 179 1288 208
rect 759 174 1288 179
rect 1288 159 1340 165
use sky130_fd_pr__nfet_g5v0d10v5_PMDTK2  sky130_fd_pr__nfet_g5v0d10v5_PMDTK2_0
timestamp 1681045192
transform 1 0 1049 0 1 776
box -108 -426 108 426
use sky130_fd_pr__nfet_g5v0d10v5_RMDT5Q  sky130_fd_pr__nfet_g5v0d10v5_RMDT5Q_0
timestamp 1681044401
transform 1 0 975 0 1 2502
box -108 -226 108 226
use sky130_fd_pr__nfet_g5v0d10v5_RMDT5Q  sky130_fd_pr__nfet_g5v0d10v5_RMDT5Q_1
timestamp 1681044401
transform 1 0 2496 0 1 2319
box -108 -226 108 226
use sky130_fd_pr__nfet_g5v0d10v5_RMDT5Q  sky130_fd_pr__nfet_g5v0d10v5_RMDT5Q_2
timestamp 1681044401
transform 1 0 2219 0 1 2315
box -108 -226 108 226
use sky130_fd_pr__nfet_g5v0d10v5_S6V9QV  sky130_fd_pr__nfet_g5v0d10v5_S6V9QV_0
timestamp 1681052864
transform 1 0 3264 0 1 909
box -345 -657 345 657
use sky130_fd_pr__nfet_g5v0d10v5_V6DT5N  sky130_fd_pr__nfet_g5v0d10v5_V6DT5N_0
timestamp 1681045192
transform 1 0 2368 0 1 1489
box -187 -226 187 226
use sky130_fd_pr__nfet_g5v0d10v5_V6DT5N  sky130_fd_pr__nfet_g5v0d10v5_V6DT5N_1
timestamp 1681045192
transform 1 0 1124 0 1 1521
box -187 -226 187 226
use sky130_fd_pr__nfet_g5v0d10v5_V6DT5N  sky130_fd_pr__nfet_g5v0d10v5_V6DT5N_2
timestamp 1681045192
transform 1 0 2525 0 1 391
box -187 -226 187 226
use sky130_fd_pr__pfet_g5v0d10v5_8FJ7Y8  sky130_fd_pr__pfet_g5v0d10v5_8FJ7Y8_0
timestamp 1681044401
transform 1 0 954 0 1 3436
box -253 -466 253 466
use sky130_fd_pr__pfet_g5v0d10v5_D4MKA2  sky130_fd_pr__pfet_g5v0d10v5_D4MKA2_0
timestamp 1681045192
transform 1 0 1499 0 1 3340
box -174 -266 174 266
use sky130_fd_pr__pfet_g5v0d10v5_D4MKA2  sky130_fd_pr__pfet_g5v0d10v5_D4MKA2_1
timestamp 1681045192
transform 1 0 1937 0 1 504
box -174 -266 174 266
use sky130_fd_pr__pfet_g5v0d10v5_D4MKA2  sky130_fd_pr__pfet_g5v0d10v5_D4MKA2_2
timestamp 1681045192
transform 1 0 1596 0 1 494
box -174 -266 174 266
use sky130_fd_pr__pfet_g5v0d10v5_D8UYD2  sky130_fd_pr__pfet_g5v0d10v5_D8UYD2_0
timestamp 1681045192
transform 1 0 1579 0 1 2607
box -253 -466 253 466
use sky130_fd_pr__pfet_g5v0d10v5_D8UYD2  sky130_fd_pr__pfet_g5v0d10v5_D8UYD2_1
timestamp 1681045192
transform 1 0 2355 0 1 3188
box -253 -466 253 466
use sky130_fd_pr__pfet_g5v0d10v5_D8UYD2  sky130_fd_pr__pfet_g5v0d10v5_D8UYD2_2
timestamp 1681045192
transform 1 0 1759 0 1 1341
box -253 -466 253 466
use sky130_fd_pr__pfet_g5v0d10v5_H9HYDU  sky130_fd_pr__pfet_g5v0d10v5_H9HYDU_0
timestamp 1681052864
transform 1 0 3259 0 1 2775
box -411 -1064 411 1102
use sky130_fd_pr__res_generic_po_RXJSZ5  sky130_fd_pr__res_generic_po_RXJSZ5_0
timestamp 1681044401
transform 1 0 313 0 1 2638
box -303 -1347 303 1347
<< labels >>
flabel metal1 s 1627 3894 1627 3894 0 FreeSans 1600 0 0 0 VDD
flabel locali s 192 971 192 971 0 FreeSans 1600 0 0 0 PLUS
flabel locali s 202 325 202 325 0 FreeSans 1600 0 0 0 VB1
flabel metal1 s 976 79 976 79 0 FreeSans 1600 0 0 0 GND
flabel metal1 s 3680 1652 3680 1652 0 FreeSans 1600 0 0 0 OUT
<< end >>
