* SPICE3 file created from opamp.ext - technology: sky130A

.subckt opamp VB1 GND VB2 PLUS VDD OUT3
X0 OUT3 a_2548_325# GND GND sky130_fd_pr__nfet_01v8 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=1
X1 a_2496_435# VB1 li_1394_1142# GND sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X2 li_604_n904# VB1 a_152_n67# GND sky130_fd_pr__nfet_01v8 ad=1.16 pd=9.16 as=0.58 ps=4.58 w=2 l=0.5
X3 a_2548_325# a_1746_n822# GND GND sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X4 GND a_1746_n822# m1_1670_n852# GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X5 m1_1412_n44# VB1 a_2548_325# VDD sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X6 li_1394_1142# VB2 GND GND sky130_fd_pr__nfet_01v8 ad=1.16 pd=9.16 as=5.22 ps=38.32 w=2 l=0.5
X7 GND VB2 li_604_n904# GND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.5
X8 m1_1670_n852# VB1 m1_875_n364# VDD sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=1.74 ps=13.16 w=2 l=0.5
X9 m1_1144_n474# OUT3 m1_875_n364# GND sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X10 m1_1412_n44# PLUS m1_1144_n474# GND sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X11 OUT3 a_2496_435# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=1
X12 m1_950_1257# GND VDD VDD sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X13 a_2496_435# a_152_n67# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=1.16 ps=8.29 w=8 l=1
X14 VDD a_152_n67# a_152_n67# VDD sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.29 as=2.32 ps=16.58 w=8 l=1
X15 GND VB2 m1_1144_n474# GND sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X16 VDD GND m1_875_n364# VDD sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X17 m1_1412_n44# GND VDD VDD sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
X18 m1_950_1257# OUT3 li_604_n904# VDD sky130_fd_pr__pfet_01v8 ad=1.74 pd=13.16 as=1.16 ps=8.58 w=4 l=1
X19 li_1394_1142# PLUS m1_950_1257# VDD sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=1
.ends
