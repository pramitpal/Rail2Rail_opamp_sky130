magic
tech sky130A
magscale 1 2
timestamp 1681046190
<< error_p >>
rect -174 1098 174 1102
rect -174 -1030 -144 1098
rect -108 1032 108 1036
rect -108 -964 -78 1032
rect 78 -964 108 1032
rect 144 -1030 174 1098
<< nwell >>
rect -144 -1064 144 1098
<< mvpmos >>
rect -50 -964 50 1036
<< mvpdiff >>
rect -108 1024 -50 1036
rect -108 -952 -96 1024
rect -62 -952 -50 1024
rect -108 -964 -50 -952
rect 50 1024 108 1036
rect 50 -952 62 1024
rect 96 -952 108 1024
rect 50 -964 108 -952
<< mvpdiffc >>
rect -96 -952 -62 1024
rect 62 -952 96 1024
<< poly >>
rect -50 1036 50 1062
rect -50 -1011 50 -964
rect -50 -1045 -34 -1011
rect 34 -1045 50 -1011
rect -50 -1061 50 -1045
<< polycont >>
rect -34 -1045 34 -1011
<< locali >>
rect -96 1024 -62 1040
rect -96 -968 -62 -952
rect 62 1024 96 1040
rect 62 -968 96 -952
rect -50 -1045 -34 -1011
rect 34 -1045 50 -1011
<< viali >>
rect -96 -952 -62 1024
rect 62 -952 96 1024
rect -34 -1045 34 -1011
<< metal1 >>
rect -102 1024 -56 1036
rect -102 -952 -96 1024
rect -62 -952 -56 1024
rect -102 -964 -56 -952
rect 56 1024 102 1036
rect 56 -952 62 1024
rect 96 -952 102 1024
rect 56 -964 102 -952
rect -46 -1011 46 -1005
rect -46 -1045 -34 -1011
rect 34 -1045 46 -1011
rect -46 -1051 46 -1045
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 10 l 0.50 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
