** sch_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/All_schematic/opamp_test/opamp.sch
.subckt opamp VOUT VINP VSSA VDDA VINN
*.PININFO VOUT:O VINP:I VSSA:B VDDA:B VINN:I
XM1 net1 net1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=8 nf=1 m=1
XM2 net2 net1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=8 nf=1 m=1
XM3 net2 net2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM4 net3 net1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=1
XM5 net6 VINN net3 VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=1
XM6 net5 VINP net3 VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=1
XM7 out net4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=8 nf=1 m=1
XM8 net4 net4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=8 nf=1 m=1
XM9 net4 Vb1 net6 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM10 out Vb1 net5 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM11 net6 net2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM12 net5 net2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM13 net7 net1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=1
XM14 net8 net1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=1
XM17 net9 net9 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM18 out2 net9 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM15 out2 Vb1 net7 VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM16 net9 Vb1 net8 VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM19 net10 net2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=1 W=4 nf=1 m=1
XM20 net8 VINN net10 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=1
XM21 net7 VINP net10 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=1
XM22 VOUT out VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=50 nf=1 m=1
XM23 VOUT out2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 nf=1 m=1
XR3 VSSA net1 VSSA sky130_fd_pr__res_generic_nd__hv W=1 L=1 mult=1 m=1
XR1 Vb1 VDDA VSSA sky130_fd_pr__res_generic_nd__hv W=1 L=1 mult=1 m=1
XR2 VSSA Vb1 VSSA sky130_fd_pr__res_generic_nd__hv W=1 L=1 mult=1 m=1
XM24 VOUT out VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=50 nf=1 m=1
XM25 VOUT out2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 nf=1 m=1
XM26 VOUT out VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=50 nf=1 m=1
XM27 VOUT out2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 nf=1 m=1
XM28 VOUT out VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=50 nf=1 m=1
XM29 VOUT out2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 nf=1 m=1
.ends
.end

.lib "/foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice.tt.red" tt


X1 VOUT VINP VSSA VDDA VOUT opamp
C1 VOUT 0 5p

V1 VSSA 0 dc 0
V2 VDDA 0 dc 3.3
******************************************************
Vin VINP 0 PWL(0 0 1u 0 1.0001u 2)

.tran 1n 10u uic

.control
set color0 = white
run

plot vinp vout xlimit 0.98u 1.05u ylimit 0 3.3
****************measuring settling_time***************
let vhi = 1.5
let vlo = 0.5
meas tran t2 WHEN v(vout)=vhi CROSS=LAST
meas tran t1 WHEN v(vout)=vlo CROSS=LAST
let slew_rate = ((vhi-vlo)/(t2-t1))/1e6
******************************************************
print slew_rate

.endc

.end
