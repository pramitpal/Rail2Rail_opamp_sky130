magic
tech sky130A
timestamp 1678605198
<< nwell >>
rect -57 -531 57 531
<< pmos >>
rect -10 -500 10 500
<< pdiff >>
rect -39 494 -10 500
rect -39 -494 -33 494
rect -16 -494 -10 494
rect -39 -500 -10 -494
rect 10 494 39 500
rect 10 -494 16 494
rect 33 -494 39 494
rect 10 -500 39 -494
<< pdiffc >>
rect -33 -494 -16 494
rect 16 -494 33 494
<< poly >>
rect -10 500 10 513
rect -10 -513 10 -500
<< locali >>
rect -33 494 -16 502
rect -33 -502 -16 -494
rect 16 494 33 502
rect 16 -502 33 -494
<< viali >>
rect -33 -494 -16 494
rect 16 -494 33 494
<< metal1 >>
rect -36 494 -13 500
rect -36 -494 -33 494
rect -16 -494 -13 494
rect -36 -500 -13 -494
rect 13 494 36 500
rect 13 -494 16 494
rect 33 -494 36 494
rect 13 -500 36 -494
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 10 l 0.2 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
