.subckt opamp
XM1 GND GND VDD VDD sky130_fd_pr__pfet_01v8 L=1000n W=3150n nf=2 m=1
XM2 net1 GND VDD VDD sky130_fd_pr__pfet_01v8 L=1000n W=3150n nf=2 m=1
XM3 net1 net1 GND GND sky130_fd_pr__nfet_01v8 L=1000n W=3150n nf=2 m=1
XM4 net2 GND VDD VDD sky130_fd_pr__pfet_01v8 L=1000n W=3150n nf=2 m=1
XM5 net6 OUT3 net2 net2 sky130_fd_pr__pfet_01v8 L=1000n W=3150n nf=2 m=1
XM6 net5 PLUS net2 net2 sky130_fd_pr__pfet_01v8 L=1000n W=3150n nf=2 m=1
XM7 net4 net3 VDD VDD sky130_fd_pr__pfet_01v8 L=1000n W=3150n nf=2 m=1
XM8 net3 net3 VDD VDD sky130_fd_pr__pfet_01v8 L=1000n W=3150n nf=2 m=1
XM9 net3 VB1 net6 net6 sky130_fd_pr__nfet_01v8 L=1000n W=3150n nf=2 m=1
XM10 net4 VB1 net5 net5 sky130_fd_pr__nfet_01v8 L=1000n W=3150n nf=2 m=1
XM11 net6 net1 GND GND sky130_fd_pr__nfet_01v8 L=1000n W=3150n nf=2 m=1
XM12 net5 net1 GND GND sky130_fd_pr__nfet_01v8 L=1000n W=3150n nf=2 m=1
XM13 net7 GND VDD VDD sky130_fd_pr__pfet_01v8 L=1000n W=3150n nf=2 m=1
XM14 net8 GND VDD VDD sky130_fd_pr__pfet_01v8 L=1000n W=3150n nf=2 m=1
XM15 net10 net10 GND GND sky130_fd_pr__nfet_01v8 L=1000n W=3150n nf=2 m=1
XM16 net9 net10 GND GND sky130_fd_pr__nfet_01v8 L=1000n W=3150n nf=2 m=1
XM17 net9 VB1 net7 net7 sky130_fd_pr__pfet_01v8 L=1000n W=3150n nf=2 m=1
XM18 net10 VB1 net8 net8 sky130_fd_pr__pfet_01v8 L=1000n W=3150n nf=2 m=1
XM19 net11 net1 GND GND sky130_fd_pr__nfet_01v8 L=1000n W=3150n nf=2 m=1
XM20 net8 OUT3 net11 net11 sky130_fd_pr__nfet_01v8 L=1000n W=3150n nf=2 m=1
XM21 net7 PLUS net11 net11 sky130_fd_pr__nfet_01v8 L=1000n W=3150n nf=2 m=1
XM22 OUT3 net4 VDD VDD sky130_fd_pr__pfet_01v8 L=1000n W=4200n nf=2 m=1
.ends
