magic
tech sky130A
magscale 1 2
timestamp 1686986091
<< error_p >>
rect -353 -466 353 466
<< nwell >>
rect -323 -462 323 462
<< mvpmos >>
rect -229 -400 -29 400
rect 29 -400 229 400
<< mvpdiff >>
rect -287 388 -229 400
rect -287 -388 -275 388
rect -241 -388 -229 388
rect -287 -400 -229 -388
rect -29 388 29 400
rect -29 -388 -17 388
rect 17 -388 29 388
rect -29 -400 29 -388
rect 229 388 287 400
rect 229 -388 241 388
rect 275 -388 287 388
rect 229 -400 287 -388
<< mvpdiffc >>
rect -275 -388 -241 388
rect -17 -388 17 388
rect 241 -388 275 388
<< poly >>
rect -229 400 -29 426
rect 29 400 229 426
rect -229 -426 -29 -400
rect 29 -426 229 -400
<< locali >>
rect -275 388 -241 404
rect -275 -404 -241 -388
rect -17 388 17 404
rect -17 -404 17 -388
rect 241 388 275 404
rect 241 -404 275 -388
<< viali >>
rect -275 -388 -241 388
rect -17 -388 17 388
rect 241 -388 275 388
<< metal1 >>
rect -281 388 -235 400
rect -281 -388 -275 388
rect -241 -388 -235 388
rect -281 -400 -235 -388
rect -23 388 23 400
rect -23 -388 -17 388
rect 17 -388 23 388
rect -23 -400 23 -388
rect 235 388 281 400
rect 235 -388 241 388
rect 275 -388 281 388
rect 235 -400 281 -388
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4 l 1 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
