magic
tech sky130A
magscale 1 2
timestamp 1681052864
<< mvnmos >>
rect -287 -831 -187 769
rect -129 -831 -29 769
rect 29 -831 129 769
rect 187 -831 287 769
<< mvndiff >>
rect -345 757 -287 769
rect -345 -819 -333 757
rect -299 -819 -287 757
rect -345 -831 -287 -819
rect -187 757 -129 769
rect -187 -819 -175 757
rect -141 -819 -129 757
rect -187 -831 -129 -819
rect -29 757 29 769
rect -29 -819 -17 757
rect 17 -819 29 757
rect -29 -831 29 -819
rect 129 757 187 769
rect 129 -819 141 757
rect 175 -819 187 757
rect 129 -831 187 -819
rect 287 757 345 769
rect 287 -819 299 757
rect 333 -819 345 757
rect 287 -831 345 -819
<< mvndiffc >>
rect -333 -819 -299 757
rect -175 -819 -141 757
rect -17 -819 17 757
rect 141 -819 175 757
rect 299 -819 333 757
<< poly >>
rect -287 841 -187 857
rect -287 807 -271 841
rect -203 807 -187 841
rect -287 769 -187 807
rect -129 841 -29 857
rect -129 807 -113 841
rect -45 807 -29 841
rect -129 769 -29 807
rect 29 841 129 857
rect 29 807 45 841
rect 113 807 129 841
rect 29 769 129 807
rect 187 841 287 857
rect 187 807 203 841
rect 271 807 287 841
rect 187 769 287 807
rect -287 -857 -187 -831
rect -129 -857 -29 -831
rect 29 -857 129 -831
rect 187 -857 287 -831
<< polycont >>
rect -271 807 -203 841
rect -113 807 -45 841
rect 45 807 113 841
rect 203 807 271 841
<< locali >>
rect -287 807 -271 841
rect -203 807 -187 841
rect -129 807 -113 841
rect -45 807 -29 841
rect 29 807 45 841
rect 113 807 129 841
rect 187 807 203 841
rect 271 807 287 841
rect -333 757 -299 773
rect -333 -835 -299 -819
rect -175 757 -141 773
rect -175 -835 -141 -819
rect -17 757 17 773
rect -17 -835 17 -819
rect 141 757 175 773
rect 141 -835 175 -819
rect 299 757 333 773
rect 299 -835 333 -819
<< viali >>
rect -271 807 -203 841
rect -113 807 -45 841
rect 45 807 113 841
rect 203 807 271 841
rect -333 -819 -299 757
rect -175 -819 -141 757
rect -17 -819 17 757
rect 141 -819 175 757
rect 299 -819 333 757
<< metal1 >>
rect -283 841 -191 847
rect -283 807 -271 841
rect -203 807 -191 841
rect -283 801 -191 807
rect -125 841 -33 847
rect -125 807 -113 841
rect -45 807 -33 841
rect -125 801 -33 807
rect 33 841 125 847
rect 33 807 45 841
rect 113 807 125 841
rect 33 801 125 807
rect 191 841 283 847
rect 191 807 203 841
rect 271 807 283 841
rect 191 801 283 807
rect -339 757 -293 769
rect -339 -819 -333 757
rect -299 -819 -293 757
rect -339 -831 -293 -819
rect -181 757 -135 769
rect -181 -819 -175 757
rect -141 -819 -135 757
rect -181 -831 -135 -819
rect -23 757 23 769
rect -23 -819 -17 757
rect 17 -819 23 757
rect -23 -831 23 -819
rect 135 757 181 769
rect 135 -819 141 757
rect 175 -819 181 757
rect 135 -831 181 -819
rect 293 757 339 769
rect 293 -819 299 757
rect 333 -819 339 757
rect 293 -831 339 -819
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 8 l 0.50 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
