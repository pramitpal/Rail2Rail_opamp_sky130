magic
tech sky130A
magscale 1 2
timestamp 1686987678
<< error_p >>
rect 36 378 252 613
rect -252 -613 -36 -378
<< mvpdiff >>
rect 102 535 186 547
rect 102 501 114 535
rect 174 501 186 535
rect 102 444 186 501
rect -186 -501 -102 -444
rect -186 -535 -174 -501
rect -114 -535 -102 -501
rect -186 -547 -102 -535
<< mvpdiffc >>
rect 114 501 174 535
rect -174 -535 -114 -501
<< mvpdiffres >>
rect -186 316 42 400
rect -186 -444 -102 316
rect -42 -316 42 316
rect 102 -316 186 444
rect -42 -400 186 -316
<< locali >>
rect 98 501 114 535
rect 174 501 190 535
rect -190 -535 -174 -501
rect -114 -535 -98 -501
<< properties >>
string gencell sky130_fd_pr__res_generic_pd__hv
string library sky130
string parameters w 0.42 l 4 m 1 nx 3 wmin 0.42 lmin 2.10 rho 197 val 6.895k dummy 0 dw 0.02 term 0.0 sterm 0.0 caplen 0.60 snake 1 guard 0 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
