* SPICE3 file created from opamp.ext - technology: sky130A

*.subckt opamp VDD VB1 GND VB2 PLUS OUT3
X0 m1_n150_n584# a_106_n270# a_2523_355# VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X1 m1_n666_n548# a_106_n270# a_130_n86# VSUBS sky130_fd_pr__nfet_01v8 ad=1.16 pd=9.16 as=0.58 ps=4.58 w=2 l=0.5
X2 a_2484_258# a_2056_n354# GND VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X3 GND a_2056_n354# a_2056_n354# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X4 a_2484_258# a_106_n270# m1_1290_528# w_1718_n12# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X5 m1_n150_n584# VB2 GND VSUBS sky130_fd_pr__nfet_01v8 ad=1.16 pd=9.16 as=4.64 ps=34.32 w=2 l=0.5
X6 GND VB2 m1_n666_n548# VSUBS sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=2 l=0.5
X7 m1_762_809# a_106_n270# a_2056_n354# w_1718_n12# sky130_fd_pr__pfet_01v8 ad=1.74 pd=13.16 as=0.58 ps=4.58 w=2 l=0.5
X8 OUT3 a_2523_355# VDD w_1718_n12# sky130_fd_pr__pfet_01v8 ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.2
X9 m1_960_n522# OUT3 m1_762_809# VSUBS sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X10 m1_1290_528# PLUS m1_960_n522# VSUBS sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X11 OUT3 a_2484_258# GND VSUBS sky130_fd_pr__nfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.2
X12 a_2523_355# a_130_n86# VDD w_n708_50# sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=1.16 ps=8.29 w=8 l=1
X13 VDD a_130_n86# a_130_n86# w_n708_50# sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.29 as=2.32 ps=16.58 w=8 l=1
X14 VDD GND m1_n406_894# w_n708_50# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X15 GND VB2 m1_960_n522# VSUBS sky130_fd_pr__nfet_01v8 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X16 m1_n406_894# OUT3 m1_n666_n548# w_n708_50# sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X17 m1_n150_n584# PLUS m1_n406_894# w_n708_50# sky130_fd_pr__pfet_01v8 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
X18 VDD GND m1_762_809# w_1718_n12# sky130_fd_pr__pfet_01v8 ad=6.96 pd=50.32 as=0 ps=0 w=4 l=1
X19 m1_1290_528# GND VDD w_1718_n12# sky130_fd_pr__pfet_01v8 ad=1.74 pd=13.16 as=0 ps=0 w=4 l=1
*.ends
