magic
tech sky130A
magscale 1 2
timestamp 1678618945
<< nwell >>
rect 0 2080 646 2081
rect 2138 2080 2504 2392
rect 0 1078 2504 2080
rect 2 506 2504 1078
rect 2 326 2174 506
rect 2 284 2170 326
rect 1524 -597 2170 284
<< psubdiff >>
rect 18 -1332 2054 -1318
rect 18 -1392 46 -1332
rect 138 -1390 448 -1332
rect 594 -1390 776 -1332
rect 138 -1392 776 -1390
rect 868 -1390 1178 -1332
rect 1324 -1390 1472 -1332
rect 868 -1392 1472 -1390
rect 1564 -1390 1874 -1332
rect 2020 -1390 2054 -1332
rect 1564 -1392 2054 -1390
rect 18 -1404 2054 -1392
<< nsubdiff >>
rect 38 1970 604 1980
rect 38 1966 426 1970
rect 38 1906 62 1966
rect 214 1910 426 1966
rect 578 1910 604 1970
rect 214 1906 604 1910
rect 38 1900 604 1906
<< psubdiffcont >>
rect 46 -1392 138 -1332
rect 448 -1390 594 -1332
rect 776 -1392 868 -1332
rect 1178 -1390 1324 -1332
rect 1472 -1392 1564 -1332
rect 1874 -1390 2020 -1332
<< nsubdiffcont >>
rect 62 1906 214 1966
rect 426 1910 578 1970
<< poly >>
rect 818 1252 878 1328
rect 726 1192 878 1252
rect 726 1178 786 1192
rect 726 1138 736 1178
rect 776 1138 786 1178
rect 726 1122 786 1138
rect 2502 489 2556 550
rect 2496 479 2562 489
rect 2496 445 2512 479
rect 2546 445 2562 479
rect 2496 435 2562 445
rect 2548 369 2614 379
rect 990 290 1080 362
rect 860 280 1080 290
rect 860 244 876 280
rect 912 244 1080 280
rect 860 234 1080 244
rect 990 174 1080 234
rect 1272 285 1362 364
rect 2548 335 2564 369
rect 2598 335 2614 369
rect 2548 325 2614 335
rect 1405 285 1471 287
rect 1272 277 1471 285
rect 1272 243 1421 277
rect 1455 243 1471 277
rect 2554 276 2608 325
rect 1272 235 1471 243
rect 1272 176 1362 235
rect 1405 233 1471 235
rect 1704 150 1772 210
rect 1970 154 2038 206
rect 1698 140 1778 150
rect 1698 92 1714 140
rect 1762 92 1778 140
rect 1698 82 1778 92
rect 1964 144 2044 154
rect 1964 96 1980 144
rect 2028 96 2044 144
rect 1964 86 2044 96
rect 162 -13 208 54
rect 438 -13 484 62
rect 152 -23 218 -13
rect 152 -57 168 -23
rect 202 -57 218 -23
rect 152 -67 218 -57
rect 428 -23 494 -13
rect 428 -57 444 -23
rect 478 -57 494 -23
rect 428 -67 494 -57
rect 118 -123 184 -113
rect 118 -157 134 -123
rect 168 -157 184 -123
rect 118 -167 184 -157
rect 478 -123 544 -113
rect 478 -157 494 -123
rect 528 -157 544 -123
rect 478 -167 544 -157
rect 128 -224 174 -167
rect 488 -226 534 -167
rect 1248 -326 1328 -316
rect 1248 -374 1264 -326
rect 1312 -374 1328 -326
rect 1248 -384 1328 -374
rect 1254 -442 1322 -384
rect 1676 -582 1744 -506
rect 1670 -592 1750 -582
rect 1980 -588 2048 -510
rect 1670 -640 1686 -592
rect 1734 -640 1750 -592
rect 1670 -650 1750 -640
rect 1974 -598 2054 -588
rect 1974 -646 1990 -598
rect 2038 -646 2054 -598
rect 1974 -656 2054 -646
rect 269 -723 335 -713
rect 269 -757 285 -723
rect 319 -757 335 -723
rect 269 -767 335 -757
rect 399 -723 465 -713
rect 399 -757 415 -723
rect 449 -757 465 -723
rect 399 -767 465 -757
rect 1748 -722 1820 -712
rect 1748 -762 1764 -722
rect 1804 -762 1820 -722
rect 282 -826 322 -767
rect 412 -826 452 -767
rect 1748 -772 1820 -762
rect 1916 -724 1988 -714
rect 1916 -764 1932 -724
rect 1972 -764 1988 -724
rect 1748 -802 1814 -772
rect 1746 -822 1814 -802
rect 1916 -804 1988 -764
rect 1916 -822 1984 -804
rect 1754 -842 1814 -822
rect 1922 -842 1982 -822
<< polycont >>
rect 736 1138 776 1178
rect 2512 445 2546 479
rect 876 244 912 280
rect 2564 335 2598 369
rect 1421 243 1455 277
rect 1714 92 1762 140
rect 1980 96 2028 144
rect 168 -57 202 -23
rect 444 -57 478 -23
rect 134 -157 168 -123
rect 494 -157 528 -123
rect 1264 -374 1312 -326
rect 1686 -640 1734 -592
rect 1990 -646 2038 -598
rect 285 -757 319 -723
rect 415 -757 449 -723
rect 1764 -762 1804 -722
rect 1932 -764 1972 -724
<< locali >>
rect 38 1972 604 1980
rect 38 1966 246 1972
rect 38 1906 62 1966
rect 214 1912 246 1966
rect 398 1970 604 1972
rect 398 1912 426 1970
rect 214 1910 426 1912
rect 578 1910 604 1970
rect 214 1906 604 1910
rect 38 1900 604 1906
rect 726 1178 786 1188
rect 720 1138 736 1178
rect 776 1138 792 1178
rect 1394 1142 1442 1240
rect 1691 1181 1929 1187
rect 1691 1139 1697 1181
rect 1739 1139 1929 1181
rect 726 668 786 1138
rect 1691 1133 1929 1139
rect 2512 489 2546 495
rect 2195 479 2556 489
rect 2195 475 2512 479
rect 676 406 920 442
rect 2195 435 2205 475
rect 2199 433 2205 435
rect 2247 445 2512 475
rect 2546 445 2556 479
rect 2247 435 2556 445
rect 2247 433 2303 435
rect 2199 427 2303 433
rect 2512 429 2546 435
rect 168 -17 202 -7
rect 444 -17 478 -7
rect 201 -23 484 -17
rect 202 -57 444 -23
rect 478 -57 484 -23
rect 201 -63 484 -57
rect 168 -73 202 -63
rect 444 -73 478 -63
rect 134 -117 168 -107
rect 494 -117 528 -107
rect 128 -123 361 -117
rect 128 -157 134 -123
rect 168 -157 361 -123
rect 128 -163 361 -157
rect 407 -123 534 -117
rect 407 -157 494 -123
rect 528 -157 534 -123
rect 407 -163 534 -157
rect 134 -173 168 -163
rect 494 -173 528 -163
rect 283 -670 336 -649
rect 283 -676 338 -670
rect 281 -684 338 -676
rect 266 -720 338 -684
rect 415 -720 449 -707
rect 266 -723 452 -720
rect 266 -757 285 -723
rect 319 -757 415 -723
rect 449 -757 452 -723
rect 266 -760 452 -757
rect 266 -770 338 -760
rect 285 -773 319 -770
rect 415 -773 449 -760
rect 676 -786 712 406
rect 2564 379 2598 385
rect 2261 369 2608 379
rect 2261 335 2564 369
rect 2598 335 2608 369
rect 2261 325 2608 335
rect 876 290 912 296
rect 872 280 922 290
rect 1421 285 1455 293
rect 872 244 876 280
rect 912 244 922 280
rect 872 234 922 244
rect 1413 277 1455 285
rect 1413 243 1421 277
rect 1413 235 1455 243
rect 876 228 912 234
rect 1421 227 1455 235
rect 1714 154 1762 156
rect 1980 154 2028 160
rect 1714 150 1830 154
rect 1704 140 1830 150
rect 1704 92 1714 140
rect 1762 92 1830 140
rect 1704 86 1830 92
rect 1898 144 2038 154
rect 1898 96 1980 144
rect 2028 96 2038 144
rect 1898 86 2038 96
rect 1704 82 1862 86
rect 1714 76 1762 82
rect 1980 80 2028 86
rect 2261 -267 2315 325
rect 2564 319 2598 325
rect 2261 -309 2267 -267
rect 2309 -309 2315 -267
rect 1264 -316 1312 -310
rect 2261 -315 2315 -309
rect 604 -822 712 -786
rect 1022 -326 1322 -316
rect 1022 -374 1264 -326
rect 1312 -374 1322 -326
rect 1022 -384 1322 -374
rect 604 -868 640 -822
rect 1022 -888 1090 -384
rect 1264 -390 1312 -384
rect 1686 -580 1734 -576
rect 1507 -582 1734 -580
rect 1507 -588 1878 -582
rect 1990 -588 2038 -582
rect 1507 -592 2048 -588
rect 1507 -640 1686 -592
rect 1734 -598 2048 -592
rect 1734 -640 1990 -598
rect 1507 -646 1990 -640
rect 2038 -646 2048 -598
rect 1507 -654 2048 -646
rect 1507 -709 1581 -654
rect 1686 -656 2048 -654
rect 1990 -662 2038 -656
rect 1764 -712 1804 -706
rect 1754 -714 1864 -712
rect 1932 -714 1972 -708
rect 1754 -722 1982 -714
rect 1754 -762 1764 -722
rect 1804 -724 1982 -722
rect 1804 -762 1932 -724
rect 1754 -764 1932 -762
rect 1972 -764 1982 -724
rect 1754 -778 1982 -764
rect 1932 -780 1972 -778
rect 812 -894 1090 -888
rect 812 -942 818 -894
rect 866 -942 1090 -894
rect 812 -948 1090 -942
rect 910 -956 1090 -948
rect 18 -1332 2062 -1316
rect 18 -1392 46 -1332
rect 138 -1334 448 -1332
rect 138 -1388 176 -1334
rect 426 -1388 448 -1334
rect 138 -1390 448 -1388
rect 594 -1390 776 -1332
rect 138 -1392 776 -1390
rect 868 -1334 1178 -1332
rect 868 -1388 906 -1334
rect 1156 -1388 1178 -1334
rect 868 -1390 1178 -1388
rect 1324 -1390 1472 -1332
rect 868 -1392 1472 -1390
rect 1564 -1334 1874 -1332
rect 1564 -1388 1602 -1334
rect 1852 -1388 1874 -1334
rect 1564 -1390 1874 -1388
rect 2020 -1390 2062 -1332
rect 1564 -1392 2062 -1390
rect 18 -1404 2062 -1392
<< viali >>
rect 246 1912 398 1972
rect 1394 1240 1442 1288
rect 1697 1139 1739 1181
rect 1929 1133 1983 1187
rect 726 608 786 668
rect 2205 433 2247 475
rect 155 -23 201 -17
rect 155 -57 168 -23
rect 168 -57 201 -23
rect 155 -63 201 -57
rect 361 -163 407 -117
rect 283 -649 336 -596
rect 816 234 872 290
rect 1455 235 1505 285
rect 1830 86 1898 154
rect 2267 -309 2309 -267
rect 604 -904 640 -868
rect 1507 -783 1581 -709
rect 818 -942 866 -894
rect 176 -1388 426 -1334
rect 906 -1388 1156 -1334
rect 1602 -1388 1852 -1334
<< metal1 >>
rect 6 1997 642 2010
rect 6 1995 688 1997
rect 6 1972 738 1995
rect 6 1912 246 1972
rect 398 1932 738 1972
rect 398 1912 642 1932
rect 6 1880 642 1912
rect 300 1652 346 1880
rect 688 1845 738 1932
rect 688 1833 1872 1845
rect 548 1751 554 1805
rect 608 1751 614 1805
rect 688 1795 2427 1833
rect 554 1642 608 1751
rect 688 1720 738 1795
rect 1822 1783 2427 1795
rect 1065 1551 1071 1605
rect 1125 1551 1131 1605
rect 1071 1415 1125 1551
rect 1071 1361 1583 1415
rect 950 1303 996 1344
rect 950 1257 1183 1303
rect 1388 1294 1448 1300
rect 1137 1111 1183 1257
rect 1382 1234 1388 1294
rect 1440 1288 1448 1294
rect 1442 1240 1448 1288
rect 1440 1234 1448 1240
rect 1388 1228 1448 1234
rect 1529 1187 1583 1361
rect 1529 1181 1751 1187
rect 1529 1139 1697 1181
rect 1739 1139 1751 1181
rect 1529 1133 1751 1139
rect 1822 1002 1872 1783
rect 1923 1187 1989 1199
rect 1923 1133 1929 1187
rect 1983 1133 2253 1187
rect 1923 1121 1989 1133
rect 714 668 798 674
rect 714 608 726 668
rect 786 608 798 668
rect 714 602 798 608
rect 726 507 786 602
rect 718 466 786 507
rect 2199 481 2253 1133
rect 2193 475 2259 481
rect 718 160 772 466
rect 2193 433 2205 475
rect 2247 433 2259 475
rect 2656 436 2704 630
rect 2193 427 2259 433
rect 2638 430 2704 436
rect 2694 374 2774 430
rect 2638 368 2704 374
rect 810 296 878 302
rect 1449 291 1511 297
rect 810 234 816 240
rect 872 234 878 240
rect 810 222 878 234
rect 1443 229 1449 291
rect 1501 285 1511 291
rect 1505 235 1511 285
rect 1501 229 1511 235
rect 1449 223 1511 229
rect 718 154 826 160
rect 45 -17 91 127
rect 149 -17 207 -5
rect 45 -63 155 -17
rect 201 -63 207 -17
rect 45 -285 91 -63
rect 149 -75 207 -63
rect 355 -111 413 -105
rect 355 -169 361 -111
rect 413 -169 419 -111
rect 355 -175 413 -169
rect 556 -252 602 113
rect 718 86 758 154
rect 718 80 826 86
rect 277 -590 342 -584
rect 277 -596 289 -590
rect 208 -714 248 -604
rect 277 -649 283 -596
rect 277 -655 289 -649
rect 342 -655 348 -590
rect 277 -661 342 -655
rect 176 -720 248 -714
rect 90 -754 248 -720
rect 395 -713 437 -567
rect 560 -630 600 -628
rect 560 -646 602 -630
rect 538 -708 604 -702
rect 496 -713 538 -710
rect 90 -756 216 -754
rect 395 -755 538 -713
rect 90 -860 126 -756
rect 76 -912 82 -860
rect 134 -912 140 -860
rect 176 -882 216 -756
rect 496 -758 538 -755
rect 498 -760 538 -758
rect 590 -760 604 -708
rect 498 -766 590 -760
rect 498 -918 538 -766
rect 598 -860 646 -856
rect 590 -912 596 -860
rect 648 -912 654 -860
rect 598 -916 646 -912
rect 330 -1300 380 -1226
rect 718 -1300 772 80
rect 1474 2 1480 5
rect 1412 -44 1480 2
rect 1474 -47 1480 -44
rect 1532 -47 1538 5
rect 1567 1 1613 295
rect 1824 160 1904 166
rect 1818 80 1824 160
rect 1892 154 1904 160
rect 1898 86 1904 154
rect 1892 80 1904 86
rect 1824 74 1904 80
rect 2085 79 2131 271
rect 2200 234 2206 286
rect 2258 234 2264 286
rect 2207 161 2257 234
rect 2656 224 2704 368
rect 2074 77 2131 79
rect 1986 5 2038 11
rect 1567 -45 1640 1
rect 1594 -107 1640 -45
rect 2074 2 2149 77
rect 2038 -11 2149 2
rect 2038 -44 2123 -11
rect 1986 -53 2038 -47
rect 2074 -116 2120 -44
rect 884 -312 930 -208
rect 875 -364 881 -312
rect 933 -364 939 -312
rect 1144 -474 1190 -192
rect 2261 -267 2315 -255
rect 1410 -312 1462 -306
rect 1498 -315 1633 -303
rect 1462 -349 1633 -315
rect 2261 -309 2267 -267
rect 2309 -309 2315 -267
rect 1462 -361 1498 -349
rect 1410 -370 1462 -364
rect 838 -558 844 -498
rect 904 -501 910 -498
rect 904 -558 921 -501
rect 844 -650 921 -558
rect 1747 -617 1797 -431
rect 847 -709 921 -650
rect 1670 -667 1797 -617
rect 1915 -645 1965 -443
rect 1501 -703 1587 -697
rect 999 -709 1073 -703
rect 847 -783 999 -709
rect 999 -789 1073 -783
rect 1495 -789 1501 -703
rect 1575 -709 1587 -703
rect 1581 -783 1587 -709
rect 1575 -789 1587 -783
rect 1501 -795 1587 -789
rect 1670 -852 1720 -667
rect 1915 -695 2040 -645
rect 1990 -724 2040 -695
rect 2261 -724 2315 -309
rect 1988 -778 2315 -724
rect 1990 -860 2040 -778
rect 812 -888 872 -882
rect 806 -948 812 -888
rect 872 -948 878 -888
rect 812 -954 872 -948
rect 1408 -1300 1452 -1224
rect 1828 -1300 1878 -1230
rect 2 -1306 2090 -1300
rect 2 -1318 2444 -1306
rect 0 -1334 2444 -1318
rect 0 -1388 176 -1334
rect 426 -1388 906 -1334
rect 1156 -1388 1602 -1334
rect 1852 -1388 2444 -1334
rect 0 -1420 2444 -1388
rect 0 -1424 2090 -1420
<< via1 >>
rect 554 1751 608 1805
rect 1071 1551 1125 1605
rect 1388 1288 1440 1294
rect 1388 1240 1394 1288
rect 1394 1240 1440 1288
rect 1388 1234 1440 1240
rect 2638 374 2694 430
rect 810 290 878 296
rect 810 240 816 290
rect 816 240 872 290
rect 872 240 878 290
rect 1449 285 1501 291
rect 1449 235 1455 285
rect 1455 235 1501 285
rect 1449 229 1501 235
rect 361 -117 413 -111
rect 361 -163 407 -117
rect 407 -163 413 -117
rect 361 -169 413 -163
rect 758 86 826 154
rect 289 -596 342 -590
rect 289 -649 336 -596
rect 336 -649 342 -596
rect 289 -655 342 -649
rect 82 -912 134 -860
rect 538 -760 590 -708
rect 596 -868 648 -860
rect 596 -904 604 -868
rect 604 -904 640 -868
rect 640 -904 648 -868
rect 596 -912 648 -904
rect 1480 -47 1532 5
rect 1824 154 1892 160
rect 1824 86 1830 154
rect 1830 86 1892 154
rect 1824 80 1892 86
rect 2206 234 2258 286
rect 1986 -47 2038 5
rect 881 -364 933 -312
rect 1410 -364 1462 -312
rect 844 -558 904 -498
rect 999 -783 1073 -709
rect 1501 -709 1575 -703
rect 1501 -783 1507 -709
rect 1507 -783 1575 -709
rect 1501 -789 1575 -783
rect 812 -894 872 -888
rect 812 -942 818 -894
rect 818 -942 866 -894
rect 866 -942 872 -894
rect 812 -948 872 -942
<< metal2 >>
rect 554 1805 608 1811
rect 608 1751 1125 1805
rect 554 1745 608 1751
rect 1071 1605 1125 1751
rect 1071 1545 1125 1551
rect 1388 1294 1440 1300
rect 638 1240 1388 1288
rect 361 -110 413 -105
rect 348 -170 357 -110
rect 417 -170 426 -110
rect 361 -175 413 -170
rect 289 -590 342 -584
rect 277 -655 286 -590
rect 346 -655 355 -590
rect 289 -661 342 -655
rect 532 -760 538 -708
rect 590 -710 596 -708
rect 638 -710 686 1240
rect 1388 1228 1440 1234
rect 816 516 2358 572
rect 816 296 872 516
rect 2302 430 2358 516
rect 2302 374 2638 430
rect 2694 374 2700 430
rect 804 240 810 296
rect 878 240 884 296
rect 1449 291 1501 297
rect 2206 286 2258 292
rect 1501 235 2206 285
rect 1449 223 1501 229
rect 2206 228 2258 234
rect 1824 160 1892 166
rect 752 86 758 154
rect 826 86 1824 154
rect 1824 74 1892 80
rect 1480 5 1532 11
rect 1980 2 1986 5
rect 1532 -44 1986 2
rect 1980 -47 1986 -44
rect 2038 -47 2044 5
rect 1480 -53 1532 -47
rect 881 -312 933 -306
rect 1404 -315 1410 -312
rect 933 -361 1410 -315
rect 1404 -364 1410 -361
rect 1462 -364 1468 -312
rect 881 -370 933 -364
rect 844 -498 904 -492
rect 837 -556 844 -500
rect 904 -556 911 -500
rect 844 -564 904 -558
rect 1501 -703 1575 -697
rect 590 -758 686 -710
rect 590 -760 596 -758
rect 993 -783 999 -709
rect 1073 -783 1501 -709
rect 1501 -795 1575 -789
rect 82 -860 134 -854
rect 596 -860 648 -854
rect 134 -904 596 -868
rect 82 -918 134 -912
rect 814 -888 870 -881
rect 596 -918 648 -912
rect 806 -948 812 -888
rect 872 -948 878 -888
rect 814 -955 870 -948
<< via2 >>
rect 357 -111 417 -110
rect 357 -169 361 -111
rect 361 -169 413 -111
rect 413 -169 417 -111
rect 357 -170 417 -169
rect 286 -655 289 -590
rect 289 -655 342 -590
rect 342 -655 346 -590
rect 846 -556 902 -500
rect 814 -946 870 -890
<< metal3 >>
rect 352 -110 422 -105
rect 352 -170 357 -110
rect 417 -170 844 -110
rect 352 -175 422 -170
rect 784 -495 844 -170
rect 784 -500 907 -495
rect 784 -556 846 -500
rect 902 -556 907 -500
rect 784 -558 907 -556
rect 841 -561 907 -558
rect 281 -590 351 -585
rect 281 -655 286 -590
rect 346 -592 351 -590
rect 346 -652 734 -592
rect 346 -655 351 -652
rect 281 -660 351 -655
rect 674 -888 734 -652
rect 809 -888 875 -885
rect 674 -890 875 -888
rect 674 -946 814 -890
rect 870 -946 875 -890
rect 674 -948 875 -946
rect 809 -951 875 -948
use sky130_fd_pr__nfet_01v8_42C9PJ  sky130_fd_pr__nfet_01v8_42C9PJ_0
timestamp 1678613396
transform 1 0 355 0 1 -1038
box -187 -226 187 226
use sky130_fd_pr__nfet_01v8_42C9PJ  sky130_fd_pr__nfet_01v8_42C9PJ_1
timestamp 1678613396
transform 1 0 1853 0 1 -1042
box -187 -226 187 226
use sky130_fd_pr__nfet_01v8_NF6LMN  sky130_fd_pr__nfet_01v8_NF6LMN_0
timestamp 1678616045
transform 1 0 2550 0 1 -744
box -158 -1026 158 1026
use sky130_fd_pr__nfet_01v8_SAC9P4  sky130_fd_pr__nfet_01v8_SAC9P4_0
timestamp 1678611711
transform 1 0 502 0 1 -438
box -108 -226 108 226
use sky130_fd_pr__nfet_01v8_SAC9P4  sky130_fd_pr__nfet_01v8_SAC9P4_1
timestamp 1678611711
transform 1 0 146 0 1 -440
box -108 -226 108 226
use sky130_fd_pr__nfet_01v8_SLJEK5  sky130_fd_pr__nfet_01v8_SLJEK5_0
timestamp 1678614268
transform 1 0 1296 0 1 -852
box -158 -426 158 426
use sky130_fd_pr__nfet_01v8_VYPHSS  sky130_fd_pr__nfet_01v8_VYPHSS_0
timestamp 1678614268
transform 1 0 1165 0 1 -38
box -287 -226 287 226
use sky130_fd_pr__pfet_01v8_7Q4LMB  sky130_fd_pr__pfet_01v8_7Q4LMB_0
timestamp 1678616045
transform 1 0 2544 0 1 1574
box -194 -1062 194 1062
use sky130_fd_pr__pfet_01v8_7Q88LS  sky130_fd_pr__pfet_01v8_7Q88LS_0
timestamp 1678614268
transform 1 0 1847 0 1 622
box -323 -462 323 462
use sky130_fd_pr__pfet_01v8_7Q88LS  sky130_fd_pr__pfet_01v8_7Q88LS_1
timestamp 1678614268
transform 1 0 1161 0 1 758
box -323 -462 323 462
use sky130_fd_pr__pfet_01v8_9Q4LM2  sky130_fd_pr__pfet_01v8_9Q4LM2_0
timestamp 1678614268
transform 1 0 844 0 1 1528
box -194 -262 194 262
use sky130_fd_pr__pfet_01v8_SK88LG  sky130_fd_pr__pfet_01v8_SK88LG_0
timestamp 1678611711
transform 1 0 323 0 1 862
box -323 -862 323 862
use sky130_fd_pr__pfet_01v8_W7GQZ7  sky130_fd_pr__pfet_01v8_W7GQZ7_0
timestamp 1678613396
transform 1 0 2018 0 1 -304
box -144 -262 144 262
use sky130_fd_pr__pfet_01v8_W7GQZ7  sky130_fd_pr__pfet_01v8_W7GQZ7_1
timestamp 1678613396
transform 1 0 1696 0 1 -298
box -144 -262 144 262
<< labels >>
flabel locali s 312 -148 312 -148 0 FreeSans 1600 0 0 0 VB1
port 1 nsew
flabel metal1 s 658 -1366 658 -1366 0 FreeSans 1600 0 0 0 GND
port 2 nsew
flabel locali s 1054 -436 1054 -436 0 FreeSans 1600 0 0 0 VB2
port 3 nsew
flabel metal1 s 2232 178 2232 178 0 FreeSans 1600 0 0 0 PLUS
port 4 nsew
flabel metal1 s 332 1902 332 1902 0 FreeSans 1600 0 0 0 VDD
port 5 nsew
flabel metal1 s 2742 398 2742 398 0 FreeSans 1600 0 0 0 OUT3
port 6 nsew
<< end >>
