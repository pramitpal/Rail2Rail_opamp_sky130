magic
tech sky130A
timestamp 1678605198
<< nwell >>
rect -97 -2531 97 2531
<< pmos >>
rect -50 -2500 50 2500
<< pdiff >>
rect -79 2494 -50 2500
rect -79 -2494 -73 2494
rect -56 -2494 -50 2494
rect -79 -2500 -50 -2494
rect 50 2494 79 2500
rect 50 -2494 56 2494
rect 73 -2494 79 2494
rect 50 -2500 79 -2494
<< pdiffc >>
rect -73 -2494 -56 2494
rect 56 -2494 73 2494
<< poly >>
rect -50 2500 50 2513
rect -50 -2513 50 -2500
<< locali >>
rect -73 2494 -56 2502
rect -73 -2502 -56 -2494
rect 56 2494 73 2502
rect 56 -2502 73 -2494
<< viali >>
rect -73 -2494 -56 2494
rect 56 -2494 73 2494
<< metal1 >>
rect -76 2494 -53 2500
rect -76 -2494 -73 2494
rect -56 -2494 -53 2494
rect -76 -2500 -53 -2494
rect 53 2494 76 2500
rect 53 -2494 56 2494
rect 73 -2494 76 2494
rect 53 -2500 76 -2494
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 50 l 1 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
