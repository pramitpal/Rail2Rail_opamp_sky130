magic
tech sky130A
magscale 1 2
timestamp 1681046190
<< error_p >>
rect -253 1598 253 1602
rect -253 -1530 -223 1598
rect -187 1532 187 1536
rect -187 -1464 -157 1532
rect 157 -1464 187 1532
rect 223 -1530 253 1598
<< nwell >>
rect -223 -1564 223 1598
<< mvpmos >>
rect -129 -1464 -29 1536
rect 29 -1464 129 1536
<< mvpdiff >>
rect -187 1524 -129 1536
rect -187 -1452 -175 1524
rect -141 -1452 -129 1524
rect -187 -1464 -129 -1452
rect -29 1524 29 1536
rect -29 -1452 -17 1524
rect 17 -1452 29 1524
rect -29 -1464 29 -1452
rect 129 1524 187 1536
rect 129 -1452 141 1524
rect 175 -1452 187 1524
rect 129 -1464 187 -1452
<< mvpdiffc >>
rect -175 -1452 -141 1524
rect -17 -1452 17 1524
rect 141 -1452 175 1524
<< poly >>
rect -129 1536 -29 1562
rect 29 1536 129 1562
rect -129 -1511 -29 -1464
rect -129 -1545 -113 -1511
rect -45 -1545 -29 -1511
rect -129 -1561 -29 -1545
rect 29 -1511 129 -1464
rect 29 -1545 45 -1511
rect 113 -1545 129 -1511
rect 29 -1561 129 -1545
<< polycont >>
rect -113 -1545 -45 -1511
rect 45 -1545 113 -1511
<< locali >>
rect -175 1524 -141 1540
rect -175 -1468 -141 -1452
rect -17 1524 17 1540
rect -17 -1468 17 -1452
rect 141 1524 175 1540
rect 141 -1468 175 -1452
rect -129 -1545 -113 -1511
rect -45 -1545 -29 -1511
rect 29 -1545 45 -1511
rect 113 -1545 129 -1511
<< viali >>
rect -175 -1452 -141 1524
rect -17 -1452 17 1524
rect 141 -1452 175 1524
rect -113 -1545 -45 -1511
rect 45 -1545 113 -1511
<< metal1 >>
rect -181 1524 -135 1536
rect -181 -1452 -175 1524
rect -141 -1452 -135 1524
rect -181 -1464 -135 -1452
rect -23 1524 23 1536
rect -23 -1452 -17 1524
rect 17 -1452 23 1524
rect -23 -1464 23 -1452
rect 135 1524 181 1536
rect 135 -1452 141 1524
rect 175 -1452 181 1524
rect 135 -1464 181 -1452
rect -125 -1511 -33 -1505
rect -125 -1545 -113 -1511
rect -45 -1545 -33 -1511
rect -125 -1551 -33 -1545
rect 33 -1511 125 -1505
rect 33 -1545 45 -1511
rect 113 -1545 125 -1511
rect 33 -1551 125 -1545
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 15 l 0.50 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
