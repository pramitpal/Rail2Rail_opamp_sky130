magic
tech sky130A
magscale 1 2
timestamp 1681053172
<< nwell >>
rect 677 3755 3685 3957
rect 697 2969 3685 3755
rect 1323 2691 3685 2969
rect 1323 2141 1832 2691
rect 1414 228 2112 1825
rect 2837 1707 3683 2691
rect 1423 226 2110 228
<< mvnmos >>
rect 925 2302 1025 2702
rect 2169 2115 2269 2515
rect 2446 2119 2546 2519
rect 995 1321 1095 1721
rect 1153 1321 1253 1721
rect 999 376 1099 1176
rect 2239 1289 2339 1689
rect 2397 1289 2497 1689
rect 2396 191 2496 591
rect 2554 191 2654 591
rect 2977 278 3077 1478
rect 3135 278 3235 1478
rect 3293 278 3393 1478
rect 3451 278 3551 1478
<< mvpmos >>
rect 825 3036 925 3836
rect 983 3036 1083 3836
rect 1449 3140 1549 3540
rect 1450 2207 1550 3007
rect 1608 2207 1708 3007
rect 2226 2788 2326 3588
rect 2384 2788 2484 3588
rect 2972 1811 3072 3811
rect 3130 1811 3230 3811
rect 3288 1811 3388 3811
rect 3446 1811 3546 3811
rect 1630 941 1730 1741
rect 1788 941 1888 1741
rect 1546 294 1646 694
rect 1887 304 1987 704
<< mvndiff >>
rect 867 2690 925 2702
rect 867 2314 879 2690
rect 913 2314 925 2690
rect 867 2302 925 2314
rect 1025 2690 1083 2702
rect 1025 2314 1037 2690
rect 1071 2314 1083 2690
rect 1025 2302 1083 2314
rect 2111 2503 2169 2515
rect 2111 2127 2123 2503
rect 2157 2127 2169 2503
rect 2111 2115 2169 2127
rect 2269 2503 2327 2515
rect 2269 2127 2281 2503
rect 2315 2127 2327 2503
rect 2269 2115 2327 2127
rect 2388 2507 2446 2519
rect 2388 2131 2400 2507
rect 2434 2131 2446 2507
rect 2388 2119 2446 2131
rect 2546 2507 2604 2519
rect 2546 2131 2558 2507
rect 2592 2131 2604 2507
rect 2546 2119 2604 2131
rect 937 1709 995 1721
rect 937 1333 949 1709
rect 983 1333 995 1709
rect 937 1321 995 1333
rect 1095 1709 1153 1721
rect 1095 1333 1107 1709
rect 1141 1333 1153 1709
rect 1095 1321 1153 1333
rect 1253 1709 1311 1721
rect 1253 1333 1265 1709
rect 1299 1333 1311 1709
rect 1253 1321 1311 1333
rect 941 1164 999 1176
rect 941 388 953 1164
rect 987 388 999 1164
rect 941 376 999 388
rect 1099 1164 1157 1176
rect 1099 388 1111 1164
rect 1145 388 1157 1164
rect 2181 1677 2239 1689
rect 2181 1301 2193 1677
rect 2227 1301 2239 1677
rect 2181 1289 2239 1301
rect 2339 1677 2397 1689
rect 2339 1301 2351 1677
rect 2385 1301 2397 1677
rect 2339 1289 2397 1301
rect 2497 1677 2555 1689
rect 2497 1301 2509 1677
rect 2543 1301 2555 1677
rect 2497 1289 2555 1301
rect 2919 1466 2977 1478
rect 1099 376 1157 388
rect 2338 579 2396 591
rect 2338 203 2350 579
rect 2384 203 2396 579
rect 2338 191 2396 203
rect 2496 579 2554 591
rect 2496 203 2508 579
rect 2542 203 2554 579
rect 2496 191 2554 203
rect 2654 579 2712 591
rect 2654 203 2666 579
rect 2700 203 2712 579
rect 2919 290 2931 1466
rect 2965 290 2977 1466
rect 2919 278 2977 290
rect 3077 1466 3135 1478
rect 3077 290 3089 1466
rect 3123 290 3135 1466
rect 3077 278 3135 290
rect 3235 1466 3293 1478
rect 3235 290 3247 1466
rect 3281 290 3293 1466
rect 3235 278 3293 290
rect 3393 1466 3451 1478
rect 3393 290 3405 1466
rect 3439 290 3451 1466
rect 3393 278 3451 290
rect 3551 1466 3609 1478
rect 3551 290 3563 1466
rect 3597 290 3609 1466
rect 3551 278 3609 290
rect 2654 191 2712 203
<< mvpdiff >>
rect 767 3824 825 3836
rect 767 3048 779 3824
rect 813 3048 825 3824
rect 767 3036 825 3048
rect 925 3824 983 3836
rect 925 3048 937 3824
rect 971 3048 983 3824
rect 925 3036 983 3048
rect 1083 3824 1141 3836
rect 1083 3048 1095 3824
rect 1129 3048 1141 3824
rect 2914 3799 2972 3811
rect 2168 3576 2226 3588
rect 1391 3528 1449 3540
rect 1391 3152 1403 3528
rect 1437 3152 1449 3528
rect 1391 3140 1449 3152
rect 1549 3528 1607 3540
rect 1549 3152 1561 3528
rect 1595 3152 1607 3528
rect 1549 3140 1607 3152
rect 1083 3036 1141 3048
rect 1392 2995 1450 3007
rect 1392 2219 1404 2995
rect 1438 2219 1450 2995
rect 1392 2207 1450 2219
rect 1550 2995 1608 3007
rect 1550 2219 1562 2995
rect 1596 2219 1608 2995
rect 1550 2207 1608 2219
rect 1708 2995 1766 3007
rect 1708 2219 1720 2995
rect 1754 2219 1766 2995
rect 2168 2800 2180 3576
rect 2214 2800 2226 3576
rect 2168 2788 2226 2800
rect 2326 3576 2384 3588
rect 2326 2800 2338 3576
rect 2372 2800 2384 3576
rect 2326 2788 2384 2800
rect 2484 3576 2542 3588
rect 2484 2800 2496 3576
rect 2530 2800 2542 3576
rect 2484 2788 2542 2800
rect 1708 2207 1766 2219
rect 2914 1823 2926 3799
rect 2960 1823 2972 3799
rect 2914 1811 2972 1823
rect 3072 3799 3130 3811
rect 3072 1823 3084 3799
rect 3118 1823 3130 3799
rect 3072 1811 3130 1823
rect 3230 3799 3288 3811
rect 3230 1823 3242 3799
rect 3276 1823 3288 3799
rect 3230 1811 3288 1823
rect 3388 3799 3446 3811
rect 3388 1823 3400 3799
rect 3434 1823 3446 3799
rect 3388 1811 3446 1823
rect 3546 3799 3604 3811
rect 3546 1823 3558 3799
rect 3592 1823 3604 3799
rect 3546 1811 3604 1823
rect 1572 1729 1630 1741
rect 1572 953 1584 1729
rect 1618 953 1630 1729
rect 1572 941 1630 953
rect 1730 1729 1788 1741
rect 1730 953 1742 1729
rect 1776 953 1788 1729
rect 1730 941 1788 953
rect 1888 1729 1946 1741
rect 1888 953 1900 1729
rect 1934 953 1946 1729
rect 1888 941 1946 953
rect 1488 682 1546 694
rect 1488 306 1500 682
rect 1534 306 1546 682
rect 1488 294 1546 306
rect 1646 682 1704 694
rect 1646 306 1658 682
rect 1692 306 1704 682
rect 1646 294 1704 306
rect 1829 692 1887 704
rect 1829 316 1841 692
rect 1875 316 1887 692
rect 1829 304 1887 316
rect 1987 692 2045 704
rect 1987 316 1999 692
rect 2033 316 2045 692
rect 1987 304 2045 316
<< mvndiffc >>
rect 879 2314 913 2690
rect 1037 2314 1071 2690
rect 2123 2127 2157 2503
rect 2281 2127 2315 2503
rect 2400 2131 2434 2507
rect 2558 2131 2592 2507
rect 949 1333 983 1709
rect 1107 1333 1141 1709
rect 1265 1333 1299 1709
rect 953 388 987 1164
rect 1111 388 1145 1164
rect 2193 1301 2227 1677
rect 2351 1301 2385 1677
rect 2509 1301 2543 1677
rect 2350 203 2384 579
rect 2508 203 2542 579
rect 2666 203 2700 579
rect 2931 290 2965 1466
rect 3089 290 3123 1466
rect 3247 290 3281 1466
rect 3405 290 3439 1466
rect 3563 290 3597 1466
<< mvpdiffc >>
rect 779 3048 813 3824
rect 937 3048 971 3824
rect 1095 3048 1129 3824
rect 1403 3152 1437 3528
rect 1561 3152 1595 3528
rect 1404 2219 1438 2995
rect 1562 2219 1596 2995
rect 1720 2219 1754 2995
rect 2180 2800 2214 3576
rect 2338 2800 2372 3576
rect 2496 2800 2530 3576
rect 2926 1823 2960 3799
rect 3084 1823 3118 3799
rect 3242 1823 3276 3799
rect 3400 1823 3434 3799
rect 3558 1823 3592 3799
rect 1584 953 1618 1729
rect 1742 953 1776 1729
rect 1900 953 1934 1729
rect 1500 306 1534 682
rect 1658 306 1692 682
rect 1841 316 1875 692
rect 1999 316 2033 692
<< psubdiff >>
rect 27 123 1213 131
rect 27 30 87 123
rect 180 30 276 123
rect 369 30 450 123
rect 543 30 633 123
rect 726 30 820 123
rect 913 30 1023 123
rect 1116 30 1213 123
rect 27 22 1213 30
<< nsubdiff >>
rect 1202 3869 1886 3877
rect 1202 3756 1243 3869
rect 1333 3756 1404 3869
rect 1517 3756 1673 3869
rect 1786 3868 1886 3869
rect 1786 3860 2734 3868
rect 1786 3768 1967 3860
rect 2059 3768 2156 3860
rect 2248 3768 2350 3860
rect 2442 3768 2555 3860
rect 2647 3768 2734 3860
rect 1786 3760 2734 3768
rect 1786 3756 1886 3760
rect 1202 3748 1886 3756
<< psubdiffcont >>
rect 87 30 180 123
rect 276 30 369 123
rect 450 30 543 123
rect 633 30 726 123
rect 820 30 913 123
rect 1023 30 1116 123
<< nsubdiffcont >>
rect 1243 3756 1333 3869
rect 1404 3756 1517 3869
rect 1673 3756 1786 3869
rect 1967 3768 2059 3860
rect 2156 3768 2248 3860
rect 2350 3768 2442 3860
rect 2555 3768 2647 3860
<< poly >>
rect 10 1341 76 1721
rect 10 1307 26 1341
rect 60 1307 76 1341
rect 10 1291 76 1307
rect 825 3836 925 3862
rect 983 3836 1083 3862
rect 2972 3811 3072 3837
rect 3130 3811 3230 3837
rect 3288 3811 3388 3837
rect 3446 3811 3546 3837
rect 2226 3588 2326 3614
rect 2384 3588 2484 3614
rect 1449 3540 1549 3566
rect 1230 3121 1284 3134
rect 1449 3121 1549 3140
rect 1230 3118 1549 3121
rect 1230 3084 1240 3118
rect 1274 3114 1549 3118
rect 1274 3084 1520 3114
rect 1230 3081 1520 3084
rect 1230 3068 1284 3081
rect 825 3010 925 3036
rect 983 3010 1083 3036
rect 716 2935 770 2950
rect 854 2935 891 3010
rect 1012 2944 1049 3010
rect 1450 3007 1550 3033
rect 1608 3007 1708 3033
rect 986 2935 1052 2944
rect 716 2934 1052 2935
rect 716 2900 726 2934
rect 760 2900 1002 2934
rect 1036 2900 1052 2934
rect 716 2898 1052 2900
rect 716 2884 770 2898
rect 986 2890 1052 2898
rect 940 2818 1006 2828
rect 940 2784 956 2818
rect 990 2784 1006 2818
rect 940 2774 1006 2784
rect 958 2732 988 2774
rect 958 2728 992 2732
rect 925 2702 1025 2728
rect 925 2276 1025 2302
rect 2226 2762 2326 2788
rect 2384 2762 2484 2788
rect 2258 2647 2304 2762
rect 2248 2643 2314 2647
rect 2421 2643 2467 2762
rect 2248 2637 2467 2643
rect 2248 2603 2264 2637
rect 2298 2603 2467 2637
rect 2248 2597 2467 2603
rect 2248 2593 2314 2597
rect 2169 2515 2269 2541
rect 2446 2519 2546 2545
rect 1450 2181 1550 2207
rect 1608 2181 1708 2207
rect 1478 2063 1518 2181
rect 1638 2064 1675 2181
rect 2169 2089 2269 2115
rect 2446 2093 2546 2119
rect 1471 2047 1525 2063
rect 1471 2013 1481 2047
rect 1515 2013 1525 2047
rect 1471 1997 1525 2013
rect 1630 2048 1684 2064
rect 1630 2014 1640 2048
rect 1674 2014 1684 2048
rect 1630 1998 1684 2014
rect 2203 2044 2246 2089
rect 2483 2044 2526 2093
rect 2203 2001 2693 2044
rect 2650 1895 2693 2001
rect 2645 1879 2699 1895
rect 1014 1845 1068 1861
rect 1014 1811 1024 1845
rect 1058 1811 1068 1845
rect 1014 1795 1068 1811
rect 1177 1841 1231 1857
rect 1177 1807 1187 1841
rect 1221 1807 1231 1841
rect 1020 1747 1062 1795
rect 1177 1791 1231 1807
rect 2337 1842 2391 1858
rect 2337 1808 2347 1842
rect 2381 1808 2391 1842
rect 2645 1845 2655 1879
rect 2689 1845 2699 1879
rect 2645 1829 2699 1845
rect 2337 1798 2391 1808
rect 1184 1747 1223 1791
rect 995 1721 1095 1747
rect 1153 1721 1253 1747
rect 1630 1741 1730 1767
rect 1788 1741 1888 1767
rect 2274 1758 2457 1798
rect 550 1341 616 1721
rect 550 1307 566 1341
rect 600 1307 616 1341
rect 550 1291 616 1307
rect 995 1295 1095 1321
rect 1153 1295 1253 1321
rect 999 1176 1099 1202
rect 2274 1715 2314 1758
rect 2417 1715 2457 1758
rect 2972 1764 3072 1811
rect 2972 1730 2988 1764
rect 3056 1730 3072 1764
rect 2239 1689 2339 1715
rect 2397 1689 2497 1715
rect 2972 1714 3072 1730
rect 3130 1764 3230 1811
rect 3130 1730 3146 1764
rect 3214 1730 3230 1764
rect 3130 1714 3230 1730
rect 3288 1764 3388 1811
rect 3288 1730 3304 1764
rect 3372 1730 3388 1764
rect 3288 1714 3388 1730
rect 3446 1764 3546 1811
rect 3446 1730 3462 1764
rect 3530 1730 3546 1764
rect 3446 1714 3546 1730
rect 2977 1550 3077 1566
rect 2977 1516 2993 1550
rect 3061 1516 3077 1550
rect 2977 1478 3077 1516
rect 3135 1550 3235 1566
rect 3135 1516 3151 1550
rect 3219 1516 3235 1550
rect 3135 1478 3235 1516
rect 3293 1550 3393 1566
rect 3293 1516 3309 1550
rect 3377 1516 3393 1550
rect 3293 1478 3393 1516
rect 3451 1550 3551 1566
rect 3451 1516 3467 1550
rect 3535 1516 3551 1550
rect 3451 1478 3551 1516
rect 2239 1263 2339 1289
rect 2397 1263 2497 1289
rect 1630 915 1730 941
rect 1788 915 1888 941
rect 1662 831 1712 915
rect 1814 831 1864 915
rect 1379 781 1864 831
rect 1379 720 1429 781
rect 2280 770 2346 778
rect 2280 768 2626 770
rect 2280 734 2296 768
rect 2330 734 2626 768
rect 2280 731 2626 734
rect 1371 710 1437 720
rect 1371 676 1387 710
rect 1421 676 1437 710
rect 1546 694 1646 720
rect 1887 704 1987 730
rect 2280 724 2346 731
rect 1371 666 1437 676
rect 999 350 1099 376
rect 1033 259 1073 350
rect 2423 617 2462 731
rect 2587 617 2626 731
rect 2396 591 2496 617
rect 2554 591 2654 617
rect 1546 268 1646 294
rect 1887 278 1987 304
rect 1026 243 1080 259
rect 1026 209 1036 243
rect 1070 209 1080 243
rect 1026 193 1080 209
rect 1351 208 1417 218
rect 1584 208 1618 268
rect 1929 208 1963 278
rect 2113 208 2179 218
rect 1351 174 1367 208
rect 1401 174 2129 208
rect 2163 174 2179 208
rect 2977 252 3077 278
rect 3135 252 3235 278
rect 3293 252 3393 278
rect 3451 252 3551 278
rect 1351 164 1417 174
rect 2113 164 2179 174
rect 2396 165 2496 191
rect 2554 165 2654 191
<< polycont >>
rect 26 1307 60 1341
rect 1240 3084 1274 3118
rect 726 2900 760 2934
rect 1002 2900 1036 2934
rect 956 2784 990 2818
rect 2264 2603 2298 2637
rect 1481 2013 1515 2047
rect 1640 2014 1674 2048
rect 1024 1811 1058 1845
rect 1187 1807 1221 1841
rect 2347 1808 2381 1842
rect 2655 1845 2689 1879
rect 566 1307 600 1341
rect 2988 1730 3056 1764
rect 3146 1730 3214 1764
rect 3304 1730 3372 1764
rect 3462 1730 3530 1764
rect 2993 1516 3061 1550
rect 3151 1516 3219 1550
rect 3309 1516 3377 1550
rect 3467 1516 3535 1550
rect 2296 734 2330 768
rect 1387 676 1421 710
rect 1036 209 1070 243
rect 1367 174 1401 208
rect 2129 174 2163 208
<< npolyres >>
rect 10 3919 184 3985
rect 10 1721 76 3919
rect 118 1891 184 3919
rect 226 3919 400 3985
rect 226 1891 292 3919
rect 118 1825 292 1891
rect 334 1891 400 3919
rect 442 3919 616 3985
rect 442 1891 508 3919
rect 334 1825 508 1891
rect 550 1721 616 3919
<< locali >>
rect 1862 3900 2788 3933
rect 1172 3869 2788 3900
rect 779 3824 813 3840
rect 775 3048 779 3088
rect 775 3032 813 3048
rect 937 3824 971 3840
rect 937 3032 971 3048
rect 1095 3824 1129 3840
rect 1172 3756 1243 3869
rect 1333 3866 1404 3869
rect 1517 3863 1673 3869
rect 1333 3756 1404 3773
rect 1517 3766 1544 3863
rect 1644 3766 1673 3863
rect 1517 3756 1673 3766
rect 1786 3862 2788 3869
rect 1786 3860 2530 3862
rect 1786 3858 1967 3860
rect 2059 3859 2156 3860
rect 1786 3765 1799 3858
rect 1876 3768 1967 3858
rect 2248 3857 2350 3860
rect 2248 3768 2271 3857
rect 2442 3770 2530 3860
rect 2651 3770 2788 3862
rect 2967 3875 3596 3923
rect 2919 3799 2967 3875
rect 2919 3783 2926 3799
rect 2442 3768 2555 3770
rect 2647 3768 2788 3770
rect 1876 3767 2036 3768
rect 2157 3767 2271 3768
rect 1876 3765 2271 3767
rect 2392 3765 2788 3768
rect 1786 3756 2788 3765
rect 1172 3718 2788 3756
rect 1862 3717 2788 3718
rect 2180 3576 2214 3592
rect 1403 3528 1437 3544
rect 1403 3136 1437 3152
rect 1561 3528 1595 3544
rect 1561 3136 1595 3152
rect 1224 3084 1237 3118
rect 1277 3084 1290 3118
rect 775 3022 812 3032
rect 725 2985 812 3022
rect 725 2950 762 2985
rect 660 2934 770 2950
rect 1002 2936 1036 2950
rect 660 2900 726 2934
rect 760 2900 776 2934
rect 660 2867 770 2900
rect 1002 2884 1036 2899
rect 660 1359 724 2867
rect 956 2818 990 2834
rect 1095 2818 1129 3048
rect 990 2784 1129 2818
rect 1404 2995 1438 3011
rect 956 2768 990 2784
rect 1038 2719 1072 2784
rect 879 2690 913 2706
rect 1037 2704 1072 2719
rect 1037 2690 1071 2704
rect 879 2298 913 2314
rect 1030 2314 1037 2509
rect 1030 2298 1071 2314
rect 1030 2146 1067 2298
rect 1404 2203 1438 2219
rect 1562 2995 1596 3011
rect 1562 2203 1596 2219
rect 1720 2995 1754 3011
rect 2171 2800 2180 2879
rect 2338 3576 2372 3592
rect 2214 2800 2217 2879
rect 2171 2643 2217 2800
rect 2338 2784 2372 2800
rect 2496 3576 2530 3592
rect 2496 2784 2530 2800
rect 2264 2643 2298 2653
rect 2171 2637 2304 2643
rect 2171 2603 2264 2637
rect 2298 2603 2304 2637
rect 2658 2606 2783 2651
rect 2670 2604 2783 2606
rect 2171 2597 2304 2603
rect 2264 2587 2298 2597
rect 2123 2503 2157 2519
rect 1754 2258 2048 2301
rect 1720 2203 1754 2219
rect 1030 2106 1918 2146
rect 1030 2076 1067 2106
rect 0 1341 110 1354
rect 0 1307 26 1341
rect 60 1307 110 1341
rect 0 1293 110 1307
rect 542 1341 724 1359
rect 542 1307 566 1341
rect 600 1307 724 1341
rect 542 1276 724 1307
rect 765 2039 1067 2076
rect 1478 2047 1518 2050
rect 1639 2048 1676 2050
rect 163 990 567 993
rect 163 956 530 990
rect 564 956 567 990
rect 163 954 567 956
rect 619 713 669 1276
rect 619 675 624 713
rect 664 675 669 713
rect 619 669 669 675
rect 185 306 682 340
rect 765 244 802 2039
rect 1465 2013 1481 2047
rect 1515 2013 1531 2047
rect 1624 2014 1640 2048
rect 1674 2014 1690 2048
rect 1478 1958 1518 2013
rect 1020 1920 1415 1958
rect 1453 1920 1518 1958
rect 1020 1918 1518 1920
rect 1020 1882 1060 1918
rect 1639 1884 1676 2014
rect 1020 1845 1062 1882
rect 1185 1845 1676 1884
rect 1878 1903 1918 2106
rect 2005 2029 2048 2258
rect 2123 2111 2157 2127
rect 2281 2503 2315 2519
rect 2281 2111 2315 2127
rect 2400 2507 2434 2523
rect 2400 2115 2434 2131
rect 2558 2507 2592 2523
rect 2736 2369 2783 2604
rect 2558 2115 2592 2131
rect 2005 2024 2560 2029
rect 2005 1990 2521 2024
rect 2555 1990 2560 2024
rect 2005 1986 2560 1990
rect 2834 1913 2883 1919
rect 2344 1903 2384 1904
rect 1878 1863 2384 1903
rect 2651 1879 2694 1884
rect 1008 1811 1024 1845
rect 1058 1811 1074 1845
rect 1185 1841 1237 1845
rect 1020 1807 1062 1811
rect 1171 1807 1187 1841
rect 1221 1807 1237 1841
rect 1185 1805 1224 1807
rect 949 1709 983 1725
rect 949 1317 983 1333
rect 1107 1709 1141 1725
rect 1107 1317 1141 1333
rect 1265 1709 1299 1725
rect 1366 1446 1405 1845
rect 2331 1842 2384 1863
rect 2639 1845 2655 1879
rect 2689 1845 2705 1879
rect 2834 1876 2840 1913
rect 2877 1876 2883 1913
rect 2331 1808 2347 1842
rect 2381 1808 2397 1842
rect 2344 1805 2384 1808
rect 1584 1729 1618 1745
rect 1265 1317 1299 1333
rect 953 1164 987 1180
rect 953 372 987 388
rect 1111 1164 1145 1180
rect 1312 853 1361 1145
rect 1584 937 1618 953
rect 1742 1729 1776 1745
rect 1742 937 1776 953
rect 1900 1729 1934 1745
rect 2193 1677 2227 1693
rect 2193 1285 2227 1301
rect 2351 1677 2385 1693
rect 2351 1285 2385 1301
rect 2509 1677 2543 1693
rect 2509 1285 2543 1301
rect 2651 1246 2694 1845
rect 2834 1676 2883 1876
rect 2960 3783 2967 3799
rect 3084 3799 3118 3815
rect 2926 1807 2960 1823
rect 3234 3799 3282 3875
rect 3548 3846 3596 3875
rect 3548 3823 3598 3846
rect 3234 3778 3242 3799
rect 3084 1807 3118 1823
rect 3276 3778 3282 3799
rect 3400 3799 3434 3815
rect 3242 1807 3276 1823
rect 3550 3799 3598 3823
rect 3550 3778 3558 3799
rect 3400 1807 3434 1823
rect 3592 3778 3598 3799
rect 3558 1807 3592 1823
rect 2972 1730 2988 1764
rect 3056 1730 3072 1764
rect 3130 1730 3146 1764
rect 3214 1730 3230 1764
rect 3288 1730 3304 1764
rect 3372 1730 3388 1764
rect 3446 1730 3462 1764
rect 3530 1730 3546 1764
rect 2834 1665 3613 1676
rect 2730 1662 3613 1665
rect 2730 1628 2733 1662
rect 2767 1628 3613 1662
rect 2730 1627 3613 1628
rect 2730 1625 2873 1627
rect 1900 937 1934 953
rect 2114 1203 2694 1246
rect 1312 846 1878 853
rect 1312 809 1835 846
rect 1872 809 1878 846
rect 1312 804 1878 809
rect 1387 718 1421 726
rect 1500 682 1534 698
rect 1387 660 1421 668
rect 1111 372 1145 388
rect 1500 290 1534 306
rect 1658 682 1692 698
rect 1658 290 1692 306
rect 1841 692 1875 708
rect 1841 300 1875 316
rect 1999 692 2033 708
rect 1999 300 2033 316
rect 876 244 1073 246
rect 765 243 1073 244
rect 765 209 1036 243
rect 1070 209 1086 243
rect 2114 226 2157 1203
rect 2208 771 2260 774
rect 2296 771 2330 784
rect 2208 768 2333 771
rect 2208 734 2296 768
rect 2330 734 2333 768
rect 2208 732 2333 734
rect 2208 594 2260 732
rect 2296 718 2330 732
rect 2807 713 2850 1520
rect 2977 1516 2993 1550
rect 3061 1516 3077 1550
rect 3135 1516 3151 1550
rect 3219 1516 3235 1550
rect 3293 1516 3309 1550
rect 3377 1516 3393 1550
rect 3451 1516 3467 1550
rect 3535 1516 3551 1550
rect 2373 708 2850 713
rect 2373 674 2377 708
rect 2411 674 2850 708
rect 2373 670 2850 674
rect 2931 1466 2965 1482
rect 2350 594 2384 595
rect 2208 579 2389 594
rect 2208 542 2350 579
rect 765 207 1073 209
rect 1367 208 1401 224
rect 876 206 1073 207
rect 1331 174 1367 208
rect 1367 158 1401 174
rect 2114 208 2186 226
rect 2114 174 2129 208
rect 2163 174 2186 208
rect 2384 542 2389 579
rect 2508 579 2542 595
rect 2350 187 2384 203
rect 2665 579 2708 670
rect 2665 535 2666 579
rect 2508 187 2542 203
rect 2700 535 2708 579
rect 2666 187 2700 203
rect 2114 164 2186 174
rect 2117 157 2186 164
rect 2805 177 2845 310
rect 3089 1466 3123 1482
rect 2931 274 2965 290
rect 3084 290 3089 322
rect 3247 1466 3281 1482
rect 3123 290 3124 322
rect 3084 177 3124 290
rect 3405 1466 3439 1482
rect 3247 274 3281 290
rect 3402 290 3405 313
rect 3563 1466 3597 1482
rect 3439 290 3442 313
rect 3402 177 3442 290
rect 3563 274 3597 290
rect 0 135 1251 157
rect 2805 137 3442 177
rect 0 131 722 135
rect 0 26 37 131
rect 141 129 543 131
rect 141 123 205 129
rect 309 123 374 129
rect 478 123 543 129
rect 647 123 722 131
rect 826 123 909 135
rect 1013 133 1251 135
rect 1013 123 1110 133
rect 180 30 205 123
rect 369 30 374 123
rect 1013 30 1023 123
rect 141 26 205 30
rect 0 24 205 26
rect 309 24 374 30
rect 478 26 543 30
rect 647 28 1110 30
rect 1214 28 1251 133
rect 647 26 1251 28
rect 478 24 1251 26
rect 0 0 1251 24
<< viali >>
rect 779 3048 813 3824
rect 937 3048 971 3824
rect 1095 3048 1129 3824
rect 1332 3773 1333 3866
rect 1333 3773 1404 3866
rect 1404 3773 1409 3866
rect 1544 3766 1644 3863
rect 2530 3860 2651 3862
rect 1799 3765 1876 3858
rect 2036 3768 2059 3859
rect 2059 3768 2156 3859
rect 2156 3768 2157 3859
rect 2271 3768 2350 3857
rect 2350 3768 2392 3857
rect 2530 3770 2555 3860
rect 2555 3770 2647 3860
rect 2647 3770 2651 3860
rect 2919 3875 2967 3923
rect 2036 3767 2157 3768
rect 2271 3765 2392 3768
rect 1403 3152 1437 3528
rect 1561 3152 1595 3528
rect 1237 3118 1277 3121
rect 1237 3084 1240 3118
rect 1240 3084 1274 3118
rect 1274 3084 1277 3118
rect 1237 3081 1277 3084
rect 1001 2934 1038 2936
rect 1001 2900 1002 2934
rect 1002 2900 1036 2934
rect 1036 2900 1038 2934
rect 1001 2899 1038 2900
rect 879 2314 913 2690
rect 1037 2314 1071 2690
rect 1404 2219 1438 2995
rect 1562 2219 1596 2995
rect 1720 2219 1754 2995
rect 2180 2800 2214 3576
rect 2338 2800 2372 3576
rect 2496 2800 2530 3576
rect 2613 2606 2658 2651
rect 110 1293 171 1354
rect 530 956 564 990
rect 624 675 664 713
rect 682 303 716 343
rect 1415 1920 1453 1958
rect 2123 2127 2157 2503
rect 2281 2127 2315 2503
rect 2400 2131 2434 2507
rect 2558 2131 2592 2507
rect 2736 2322 2783 2369
rect 2521 1990 2555 2024
rect 949 1333 983 1709
rect 1107 1333 1141 1709
rect 1265 1333 1299 1709
rect 2840 1876 2877 1913
rect 1366 1407 1405 1446
rect 953 388 987 1164
rect 1111 388 1145 1164
rect 1312 1145 1361 1194
rect 1584 953 1618 1729
rect 1742 953 1776 1729
rect 1900 953 1934 1729
rect 2193 1301 2227 1677
rect 2351 1301 2385 1677
rect 2509 1301 2543 1677
rect 2926 1823 2960 3799
rect 3084 1823 3118 3799
rect 3242 1823 3276 3799
rect 3400 1823 3434 3799
rect 3558 1823 3592 3799
rect 2988 1730 3056 1764
rect 3146 1730 3214 1764
rect 3304 1730 3372 1764
rect 3462 1730 3530 1764
rect 2733 1628 2767 1662
rect 3613 1627 3662 1676
rect 2807 1520 2850 1563
rect 1835 809 1872 846
rect 1379 710 1429 718
rect 1379 676 1387 710
rect 1387 676 1421 710
rect 1421 676 1429 710
rect 1379 668 1429 676
rect 1500 306 1534 682
rect 1658 306 1692 682
rect 1841 316 1875 692
rect 1999 316 2033 692
rect 2993 1516 3061 1550
rect 3151 1516 3219 1550
rect 3309 1516 3377 1550
rect 3467 1516 3535 1550
rect 2377 674 2411 708
rect 1297 174 1331 208
rect 2350 203 2384 579
rect 2508 203 2542 579
rect 2666 203 2700 579
rect 2805 310 2845 350
rect 2931 290 2965 1466
rect 3089 290 3123 1466
rect 3247 290 3281 1466
rect 3405 290 3439 1466
rect 3563 290 3597 1466
rect 37 123 141 131
rect 205 123 309 129
rect 374 123 478 129
rect 543 123 647 131
rect 722 123 826 135
rect 909 123 1013 135
rect 1110 123 1214 133
rect 37 30 87 123
rect 87 30 141 123
rect 205 30 276 123
rect 276 30 309 123
rect 374 30 450 123
rect 450 30 478 123
rect 543 30 633 123
rect 633 30 647 123
rect 722 30 726 123
rect 726 30 820 123
rect 820 30 826 123
rect 909 30 913 123
rect 913 30 1013 123
rect 1110 30 1116 123
rect 1116 30 1214 123
rect 37 26 141 30
rect 205 24 309 30
rect 374 24 478 30
rect 543 26 647 30
rect 1110 28 1214 30
<< metal1 >>
rect 1862 3932 2788 3933
rect 931 3923 2788 3932
rect 2913 3923 2973 3935
rect 931 3885 2919 3923
rect 773 3824 819 3836
rect 773 3048 779 3824
rect 813 3048 819 3824
rect 773 3036 819 3048
rect 931 3824 978 3885
rect 1166 3875 2919 3885
rect 2967 3875 2973 3923
rect 1166 3866 2788 3875
rect 931 3048 937 3824
rect 971 3811 978 3824
rect 1089 3824 1135 3836
rect 971 3048 977 3811
rect 931 3036 977 3048
rect 1089 3048 1095 3824
rect 1129 3048 1135 3824
rect 1166 3773 1332 3866
rect 1409 3863 2788 3866
rect 2913 3863 2973 3875
rect 3068 3872 3074 3924
rect 3126 3875 3445 3924
rect 3126 3872 3132 3875
rect 1409 3773 1544 3863
rect 1166 3766 1544 3773
rect 1644 3862 2788 3863
rect 1644 3859 2530 3862
rect 1644 3858 2036 3859
rect 1644 3766 1799 3858
rect 1166 3765 1799 3766
rect 1876 3767 2036 3858
rect 2157 3857 2530 3859
rect 2157 3767 2271 3857
rect 1876 3765 2271 3767
rect 2392 3770 2530 3857
rect 2651 3770 2788 3862
rect 2392 3765 2788 3770
rect 1166 3718 2788 3765
rect 1390 3528 1443 3718
rect 1862 3717 2788 3718
rect 2920 3799 2966 3811
rect 1390 3522 1403 3528
rect 1397 3152 1403 3522
rect 1437 3152 1443 3528
rect 1397 3140 1443 3152
rect 1555 3528 1601 3540
rect 1555 3152 1561 3528
rect 1595 3165 1601 3528
rect 1595 3152 1605 3165
rect 1555 3140 1605 3152
rect 1225 3121 1289 3127
rect 1225 3081 1237 3121
rect 1277 3081 1289 3121
rect 1225 3075 1289 3081
rect 1089 3036 1135 3048
rect 995 2937 1044 2948
rect 1237 2937 1277 3075
rect 1557 3007 1605 3140
rect 995 2936 1277 2937
rect 995 2899 1001 2936
rect 1038 2900 1277 2936
rect 1398 2995 1444 3007
rect 1038 2899 1044 2900
rect 995 2887 1044 2899
rect 873 2690 919 2702
rect 873 2396 879 2690
rect 861 2314 879 2396
rect 913 2396 919 2690
rect 1031 2690 1077 2702
rect 913 2314 922 2396
rect 861 2171 922 2314
rect 1031 2314 1037 2690
rect 1071 2314 1077 2690
rect 1031 2302 1077 2314
rect 1398 2257 1404 2995
rect 745 2117 922 2171
rect 1383 2219 1404 2257
rect 1438 2219 1444 2995
rect 1383 2207 1444 2219
rect 1556 2995 1605 3007
rect 1556 2219 1562 2995
rect 1596 2989 1605 2995
rect 1714 2995 1760 3007
rect 1596 2219 1602 2989
rect 1556 2207 1602 2219
rect 1714 2219 1720 2995
rect 1754 2219 1760 2995
rect 1866 2399 1910 3717
rect 2174 3576 2220 3588
rect 2174 2800 2180 3576
rect 2214 2800 2220 3576
rect 2331 3576 2378 3717
rect 2826 3620 2832 3672
rect 2884 3620 2890 3672
rect 2331 3541 2338 3576
rect 2174 2788 2220 2800
rect 2332 2800 2338 3541
rect 2372 2800 2378 3576
rect 2332 2788 2378 2800
rect 2490 3576 2536 3588
rect 2490 2800 2496 3576
rect 2530 2831 2536 3576
rect 2530 2800 2550 2831
rect 2490 2788 2550 2800
rect 2174 2676 2219 2788
rect 2174 2631 2322 2676
rect 2277 2515 2322 2631
rect 2505 2652 2550 2788
rect 2607 2652 2664 2663
rect 2505 2651 2664 2652
rect 2505 2627 2613 2651
rect 2117 2503 2163 2515
rect 1856 2347 1862 2399
rect 1914 2347 1920 2399
rect 1714 2207 1760 2219
rect 745 2110 921 2117
rect 745 1628 806 2110
rect 1383 2084 1426 2207
rect 2117 2127 2123 2503
rect 2157 2127 2163 2503
rect 2117 2115 2163 2127
rect 2275 2503 2322 2515
rect 2275 2127 2281 2503
rect 2315 2483 2322 2503
rect 2392 2607 2613 2627
rect 2392 2582 2550 2607
rect 2607 2606 2613 2607
rect 2658 2606 2664 2651
rect 2607 2594 2664 2606
rect 2392 2519 2437 2582
rect 2392 2507 2440 2519
rect 2392 2484 2400 2507
rect 2315 2127 2321 2483
rect 2275 2115 2321 2127
rect 2394 2131 2400 2484
rect 2434 2131 2440 2507
rect 2394 2119 2440 2131
rect 2552 2507 2598 2519
rect 2552 2131 2558 2507
rect 2592 2154 2598 2507
rect 2724 2369 2795 2375
rect 2724 2322 2736 2369
rect 2783 2322 2795 2369
rect 2724 2316 2795 2322
rect 2592 2131 2600 2154
rect 2552 2119 2600 2131
rect 1383 2078 1897 2084
rect 1383 2041 2048 2078
rect 1789 2040 2048 2041
rect 2118 2040 2161 2115
rect 1789 2035 2235 2040
rect 2005 1997 2235 2035
rect 2557 2030 2600 2119
rect 1784 1983 1836 1989
rect 1403 1958 1465 1964
rect 1403 1920 1415 1958
rect 1453 1920 1465 1958
rect 1403 1914 1465 1920
rect 1740 1931 1784 1936
rect 1740 1925 1836 1931
rect 412 1567 806 1628
rect 943 1709 989 1721
rect 104 1355 177 1366
rect 412 1355 473 1567
rect 835 1454 887 1460
rect 670 1409 835 1448
rect 104 1354 479 1355
rect 104 1293 110 1354
rect 171 1339 479 1354
rect 171 1294 481 1339
rect 171 1293 177 1294
rect 104 1281 177 1293
rect 435 157 481 1294
rect 518 992 576 996
rect 670 992 709 1409
rect 835 1396 887 1402
rect 943 1376 949 1709
rect 937 1333 949 1376
rect 983 1333 989 1709
rect 937 1321 989 1333
rect 1101 1709 1147 1721
rect 1101 1333 1107 1709
rect 1141 1356 1147 1709
rect 1259 1709 1305 1721
rect 1141 1333 1154 1356
rect 1101 1321 1154 1333
rect 937 1282 986 1321
rect 842 1233 986 1282
rect 842 1193 891 1233
rect 834 1141 840 1193
rect 892 1141 898 1193
rect 1106 1176 1154 1321
rect 1259 1333 1265 1709
rect 1299 1333 1305 1709
rect 1409 1624 1459 1914
rect 1740 1892 1832 1925
rect 1740 1741 1784 1892
rect 1578 1729 1624 1741
rect 1402 1572 1408 1624
rect 1460 1572 1466 1624
rect 1360 1453 1411 1458
rect 1354 1401 1360 1453
rect 1412 1401 1418 1453
rect 1360 1395 1411 1401
rect 1259 1277 1305 1333
rect 1259 1231 1364 1277
rect 1312 1200 1361 1231
rect 947 1164 993 1176
rect 518 990 709 992
rect 518 956 530 990
rect 564 956 709 990
rect 518 953 709 956
rect 518 950 576 953
rect 618 719 670 725
rect 612 667 618 719
rect 670 667 676 719
rect 618 663 670 667
rect 947 388 953 1164
rect 987 388 993 1164
rect 676 349 728 355
rect 670 297 676 349
rect 676 291 728 297
rect 947 157 993 388
rect 1105 1164 1154 1176
rect 1105 388 1111 1164
rect 1145 1158 1154 1164
rect 1300 1194 1373 1200
rect 1145 388 1151 1158
rect 1300 1145 1312 1194
rect 1361 1145 1373 1194
rect 1300 1139 1373 1145
rect 1578 986 1584 1729
rect 1576 953 1584 986
rect 1618 986 1624 1729
rect 1736 1729 1784 1741
rect 1618 953 1625 986
rect 1285 917 1337 923
rect 1576 915 1625 953
rect 1736 953 1742 1729
rect 1776 1712 1784 1729
rect 1894 1729 1940 1741
rect 1776 953 1782 1712
rect 1894 965 1900 1729
rect 1736 941 1782 953
rect 1892 953 1900 965
rect 1934 965 1940 1729
rect 2192 1689 2235 1997
rect 2509 2024 2600 2030
rect 2509 1990 2521 2024
rect 2555 1990 2600 2024
rect 2509 1985 2600 1990
rect 2509 1984 2567 1985
rect 2512 1689 2555 1984
rect 2736 1773 2783 2316
rect 2834 1913 2883 3620
rect 2834 1876 2840 1913
rect 2877 1876 2883 1913
rect 2834 1864 2883 1876
rect 2920 1823 2926 3799
rect 2960 1823 2966 3799
rect 3075 3799 3124 3872
rect 3075 3796 3084 3799
rect 2920 1811 2966 1823
rect 3078 1823 3084 3796
rect 3118 1823 3124 3799
rect 3078 1811 3124 1823
rect 3236 3799 3282 3811
rect 3392 3800 3441 3875
rect 3236 1823 3242 3799
rect 3276 1823 3282 3799
rect 3236 1811 3282 1823
rect 3394 3799 3440 3800
rect 3394 1823 3400 3799
rect 3434 1823 3440 3799
rect 3394 1811 3440 1823
rect 3552 3799 3598 3811
rect 3552 1823 3558 3799
rect 3592 1823 3598 3799
rect 3552 1811 3598 1823
rect 2736 1764 3542 1773
rect 2736 1730 2988 1764
rect 3056 1730 3146 1764
rect 3214 1730 3304 1764
rect 3372 1730 3462 1764
rect 3530 1730 3542 1764
rect 2736 1726 3542 1730
rect 2951 1718 3542 1726
rect 2187 1677 2235 1689
rect 2187 1301 2193 1677
rect 2227 1645 2235 1677
rect 2345 1677 2391 1689
rect 2227 1301 2233 1645
rect 2345 1307 2351 1677
rect 2187 1289 2233 1301
rect 2343 1301 2351 1307
rect 2385 1307 2391 1677
rect 2503 1677 2555 1689
rect 2385 1301 2393 1307
rect 2343 1063 2393 1301
rect 2503 1301 2509 1677
rect 2543 1654 2555 1677
rect 3574 1676 3699 1703
rect 2721 1662 2779 1668
rect 2543 1301 2549 1654
rect 2582 1624 2634 1630
rect 2721 1628 2733 1662
rect 2767 1628 2779 1662
rect 2721 1623 2779 1628
rect 2634 1622 2779 1623
rect 3574 1627 3613 1676
rect 3662 1627 3699 1676
rect 2634 1573 2770 1622
rect 3574 1596 3699 1627
rect 2582 1566 2634 1572
rect 2503 1289 2549 1301
rect 2730 1340 2770 1573
rect 2801 1563 2856 1575
rect 2970 1563 3561 1565
rect 2801 1520 2807 1563
rect 2850 1550 3561 1563
rect 2850 1520 2993 1550
rect 2801 1508 2856 1520
rect 2970 1516 2993 1520
rect 3061 1516 3151 1550
rect 3219 1516 3309 1550
rect 3377 1516 3467 1550
rect 3535 1516 3561 1550
rect 2970 1510 3561 1516
rect 2925 1466 2971 1478
rect 2730 1300 2845 1340
rect 2343 1013 2551 1063
rect 2343 1009 2393 1013
rect 1934 953 1941 965
rect 1337 866 1625 915
rect 1285 859 1337 865
rect 1576 846 1625 866
rect 1892 852 1941 953
rect 1823 846 1941 852
rect 1576 797 1702 846
rect 1823 809 1835 846
rect 1872 809 1941 846
rect 1823 803 1941 809
rect 1373 724 1435 730
rect 1367 662 1373 724
rect 1425 718 1435 724
rect 1429 668 1435 718
rect 1653 694 1702 797
rect 1425 662 1435 668
rect 1373 656 1435 662
rect 1494 682 1540 694
rect 1105 376 1151 388
rect 1494 306 1500 682
rect 1534 306 1540 682
rect 1494 294 1540 306
rect 1652 682 1702 694
rect 1829 704 1878 803
rect 2365 712 2423 714
rect 2216 708 2423 712
rect 1829 692 1881 704
rect 1829 684 1841 692
rect 1652 306 1658 682
rect 1692 676 1702 682
rect 1692 306 1698 676
rect 1652 294 1698 306
rect 1835 316 1841 684
rect 1875 316 1881 692
rect 1835 304 1881 316
rect 1993 692 2039 704
rect 1993 316 1999 692
rect 2033 338 2039 692
rect 2216 674 2377 708
rect 2411 674 2423 708
rect 2216 669 2423 674
rect 2033 316 2072 338
rect 1993 304 2072 316
rect 1291 217 1337 220
rect 1282 165 1288 217
rect 1340 165 1346 217
rect 1291 162 1337 165
rect 0 135 1251 157
rect 0 131 722 135
rect 0 26 37 131
rect 141 129 543 131
rect 141 26 205 129
rect 0 24 205 26
rect 309 24 374 129
rect 478 26 543 129
rect 647 30 722 131
rect 826 30 909 135
rect 1013 133 1251 135
rect 1013 30 1110 133
rect 647 28 1110 30
rect 1214 129 1251 133
rect 1494 150 1532 294
rect 1996 290 2072 304
rect 2216 290 2259 669
rect 2365 668 2423 669
rect 1996 247 2259 290
rect 2344 579 2390 591
rect 2344 203 2350 579
rect 2384 203 2390 579
rect 2501 579 2551 1013
rect 2501 538 2508 579
rect 2344 191 2390 203
rect 2502 203 2508 538
rect 2542 538 2551 579
rect 2660 579 2706 591
rect 2542 256 2548 538
rect 2542 203 2553 256
rect 2502 191 2553 203
rect 2660 203 2666 579
rect 2700 203 2706 579
rect 2805 356 2845 1300
rect 2793 350 2857 356
rect 2793 310 2805 350
rect 2845 310 2857 350
rect 2793 304 2857 310
rect 2925 290 2931 1466
rect 2965 290 2971 1466
rect 2925 287 2971 290
rect 3083 1466 3129 1478
rect 3083 290 3089 1466
rect 3123 290 3129 1466
rect 2925 286 2972 287
rect 2925 255 2978 286
rect 3083 278 3129 290
rect 3241 1466 3287 1478
rect 3241 290 3247 1466
rect 3281 320 3287 1466
rect 3399 1466 3445 1478
rect 3281 290 3292 320
rect 3241 278 3292 290
rect 3399 290 3405 1466
rect 3439 290 3445 1466
rect 3399 278 3445 290
rect 3557 1466 3603 1478
rect 3557 290 3563 1466
rect 3597 335 3603 1466
rect 3597 290 3607 335
rect 3557 278 3607 290
rect 2660 191 2706 203
rect 2932 201 2978 255
rect 3246 201 3292 278
rect 3561 201 3607 278
rect 2348 150 2386 191
rect 1214 75 1260 129
rect 1494 112 2386 150
rect 2507 75 2553 191
rect 2932 155 3607 201
rect 2932 75 2978 155
rect 1214 29 2978 75
rect 1214 28 1260 29
rect 647 26 1260 28
rect 478 24 1260 26
rect 0 0 1260 24
<< via1 >>
rect 3074 3872 3126 3924
rect 2832 3620 2884 3672
rect 1862 2347 1914 2399
rect 1784 1931 1836 1983
rect 835 1402 887 1454
rect 840 1141 892 1193
rect 1408 1572 1460 1624
rect 1360 1446 1412 1453
rect 1360 1407 1366 1446
rect 1366 1407 1405 1446
rect 1405 1407 1412 1446
rect 1360 1401 1412 1407
rect 618 713 670 719
rect 618 675 624 713
rect 624 675 664 713
rect 664 675 670 713
rect 618 667 670 675
rect 676 343 728 349
rect 676 303 682 343
rect 682 303 716 343
rect 716 303 728 343
rect 676 297 728 303
rect 1285 865 1337 917
rect 2582 1572 2634 1624
rect 1373 718 1425 724
rect 1373 668 1379 718
rect 1379 668 1425 718
rect 1373 662 1425 668
rect 1288 208 1340 217
rect 1288 174 1297 208
rect 1297 174 1331 208
rect 1331 174 1340 208
rect 1288 165 1340 174
<< metal2 >>
rect 3074 3924 3126 3930
rect 2833 3874 3074 3923
rect 2833 3678 2882 3874
rect 3074 3866 3126 3872
rect 2832 3672 2884 3678
rect 2832 3614 2884 3620
rect 1862 2399 1914 2405
rect 1788 2351 1862 2395
rect 1788 1983 1832 2351
rect 1862 2341 1914 2347
rect 1778 1931 1784 1983
rect 1836 1931 1842 1983
rect 1408 1624 1460 1630
rect 1405 1573 1408 1623
rect 2576 1623 2582 1624
rect 1460 1573 2582 1623
rect 2576 1572 2582 1573
rect 2634 1572 2640 1624
rect 1408 1566 1460 1572
rect 829 1402 835 1454
rect 887 1447 893 1454
rect 1360 1453 1412 1459
rect 887 1408 1360 1447
rect 887 1402 893 1408
rect 1360 1395 1412 1401
rect 840 1193 892 1199
rect 892 1189 1328 1191
rect 892 1142 1336 1189
rect 840 1135 892 1141
rect 1287 917 1336 1142
rect 1279 865 1285 917
rect 1337 865 1343 917
rect 618 719 670 725
rect 1373 724 1425 730
rect 670 668 1373 718
rect 618 661 670 667
rect 1373 656 1425 662
rect 670 297 676 349
rect 728 297 734 349
rect 685 208 719 297
rect 1288 217 1340 223
rect 685 179 1288 208
rect 759 174 1288 179
rect 1288 159 1340 165
<< labels >>
flabel metal1 s 1627 3894 1627 3894 0 FreeSans 1600 0 0 0 VDD
port 1 nsew
flabel locali s 192 971 192 971 0 FreeSans 1600 0 0 0 PLUS
port 2 nsew
flabel locali s 202 325 202 325 0 FreeSans 1600 0 0 0 VB1
port 3 nsew
flabel metal1 s 976 79 976 79 0 FreeSans 1600 0 0 0 GND
port 4 nsew
flabel metal1 s 3680 1652 3680 1652 0 FreeSans 1600 0 0 0 OUT
port 5 nsew
<< end >>
