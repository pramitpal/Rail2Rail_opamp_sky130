magic
tech sky130A
magscale 1 2
timestamp 1686987678
<< xpolycontact >>
rect 131 154 201 586
rect -201 -586 -131 -154
<< xpolyres >>
rect -201 20 35 50
rect 131 20 201 154
rect -201 -20 201 20
rect -201 -154 -131 -20
rect -35 -50 201 -20
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p35
string library sky130
string parameters w 0.35 l 0.5 m 1 nx 3 wmin 0.350 lmin 0.50 rho 2000 val 13.646k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.350 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 1 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
