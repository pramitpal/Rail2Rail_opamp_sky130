magic
tech sky130A
magscale 1 2
timestamp 1681052864
<< mvnmos >>
rect -287 -631 -187 569
rect -129 -631 -29 569
rect 29 -631 129 569
rect 187 -631 287 569
<< mvndiff >>
rect -345 557 -287 569
rect -345 -619 -333 557
rect -299 -619 -287 557
rect -345 -631 -287 -619
rect -187 557 -129 569
rect -187 -619 -175 557
rect -141 -619 -129 557
rect -187 -631 -129 -619
rect -29 557 29 569
rect -29 -619 -17 557
rect 17 -619 29 557
rect -29 -631 29 -619
rect 129 557 187 569
rect 129 -619 141 557
rect 175 -619 187 557
rect 129 -631 187 -619
rect 287 557 345 569
rect 287 -619 299 557
rect 333 -619 345 557
rect 287 -631 345 -619
<< mvndiffc >>
rect -333 -619 -299 557
rect -175 -619 -141 557
rect -17 -619 17 557
rect 141 -619 175 557
rect 299 -619 333 557
<< poly >>
rect -287 641 -187 657
rect -287 607 -271 641
rect -203 607 -187 641
rect -287 569 -187 607
rect -129 641 -29 657
rect -129 607 -113 641
rect -45 607 -29 641
rect -129 569 -29 607
rect 29 641 129 657
rect 29 607 45 641
rect 113 607 129 641
rect 29 569 129 607
rect 187 641 287 657
rect 187 607 203 641
rect 271 607 287 641
rect 187 569 287 607
rect -287 -657 -187 -631
rect -129 -657 -29 -631
rect 29 -657 129 -631
rect 187 -657 287 -631
<< polycont >>
rect -271 607 -203 641
rect -113 607 -45 641
rect 45 607 113 641
rect 203 607 271 641
<< locali >>
rect -287 607 -271 641
rect -203 607 -187 641
rect -129 607 -113 641
rect -45 607 -29 641
rect 29 607 45 641
rect 113 607 129 641
rect 187 607 203 641
rect 271 607 287 641
rect -333 557 -299 573
rect -333 -635 -299 -619
rect -175 557 -141 573
rect -175 -635 -141 -619
rect -17 557 17 573
rect -17 -635 17 -619
rect 141 557 175 573
rect 141 -635 175 -619
rect 299 557 333 573
rect 299 -635 333 -619
<< viali >>
rect -271 607 -203 641
rect -113 607 -45 641
rect 45 607 113 641
rect 203 607 271 641
rect -333 -619 -299 557
rect -175 -619 -141 557
rect -17 -619 17 557
rect 141 -619 175 557
rect 299 -619 333 557
<< metal1 >>
rect -283 641 -191 647
rect -283 607 -271 641
rect -203 607 -191 641
rect -283 601 -191 607
rect -125 641 -33 647
rect -125 607 -113 641
rect -45 607 -33 641
rect -125 601 -33 607
rect 33 641 125 647
rect 33 607 45 641
rect 113 607 125 641
rect 33 601 125 607
rect 191 641 283 647
rect 191 607 203 641
rect 271 607 283 641
rect 191 601 283 607
rect -339 557 -293 569
rect -339 -619 -333 557
rect -299 -619 -293 557
rect -339 -631 -293 -619
rect -181 557 -135 569
rect -181 -619 -175 557
rect -141 -619 -135 557
rect -181 -631 -135 -619
rect -23 557 23 569
rect -23 -619 -17 557
rect 17 -619 23 557
rect -23 -631 23 -619
rect 135 557 181 569
rect 135 -619 141 557
rect 175 -619 181 557
rect 135 -631 181 -619
rect 293 557 339 569
rect 293 -619 299 557
rect 333 -619 339 557
rect 293 -631 339 -619
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 6 l 0.50 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
