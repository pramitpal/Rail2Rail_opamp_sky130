magic
tech sky130A
timestamp 1686980626
<< error_p >>
rect -370 -433 370 433
<< nwell >>
rect -355 -431 355 431
<< mvpmos >>
rect -308 -400 -208 400
rect -179 -400 -79 400
rect -50 -400 50 400
rect 79 -400 179 400
rect 208 -400 308 400
<< mvpdiff >>
rect -337 394 -308 400
rect -337 -394 -331 394
rect -314 -394 -308 394
rect -337 -400 -308 -394
rect -208 394 -179 400
rect -208 -394 -202 394
rect -185 -394 -179 394
rect -208 -400 -179 -394
rect -79 394 -50 400
rect -79 -394 -73 394
rect -56 -394 -50 394
rect -79 -400 -50 -394
rect 50 394 79 400
rect 50 -394 56 394
rect 73 -394 79 394
rect 50 -400 79 -394
rect 179 394 208 400
rect 179 -394 185 394
rect 202 -394 208 394
rect 179 -400 208 -394
rect 308 394 337 400
rect 308 -394 314 394
rect 331 -394 337 394
rect 308 -400 337 -394
<< mvpdiffc >>
rect -331 -394 -314 394
rect -202 -394 -185 394
rect -73 -394 -56 394
rect 56 -394 73 394
rect 185 -394 202 394
rect 314 -394 331 394
<< poly >>
rect -308 400 -208 413
rect -179 400 -79 413
rect -50 400 50 413
rect 79 400 179 413
rect 208 400 308 413
rect -308 -413 -208 -400
rect -179 -413 -79 -400
rect -50 -413 50 -400
rect 79 -413 179 -400
rect 208 -413 308 -400
<< locali >>
rect -331 394 -314 402
rect -331 -402 -314 -394
rect -202 394 -185 402
rect -202 -402 -185 -394
rect -73 394 -56 402
rect -73 -402 -56 -394
rect 56 394 73 402
rect 56 -402 73 -394
rect 185 394 202 402
rect 185 -402 202 -394
rect 314 394 331 402
rect 314 -402 331 -394
<< viali >>
rect -331 -394 -314 394
rect -202 -394 -185 394
rect -73 -394 -56 394
rect 56 -394 73 394
rect 185 -394 202 394
rect 314 -394 331 394
<< metal1 >>
rect -334 394 -311 400
rect -334 -394 -331 394
rect -314 -394 -311 394
rect -334 -400 -311 -394
rect -205 394 -182 400
rect -205 -394 -202 394
rect -185 -394 -182 394
rect -205 -400 -182 -394
rect -76 394 -53 400
rect -76 -394 -73 394
rect -56 -394 -53 394
rect -76 -400 -53 -394
rect 53 394 76 400
rect 53 -394 56 394
rect 73 -394 76 394
rect 53 -400 76 -394
rect 182 394 205 400
rect 182 -394 185 394
rect 202 -394 205 394
rect 182 -400 205 -394
rect 311 394 334 400
rect 311 -394 314 394
rect 331 -394 334 394
rect 311 -400 334 -394
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 8 l 1 m 1 nf 5 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
