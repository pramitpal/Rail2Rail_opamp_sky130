magic
tech sky130A
magscale 1 2
timestamp 1678601982
<< nwell >>
rect -323 -862 323 862
<< pmos >>
rect -229 -800 -29 800
rect 29 -800 229 800
<< pdiff >>
rect -287 788 -229 800
rect -287 -788 -275 788
rect -241 -788 -229 788
rect -287 -800 -229 -788
rect -29 788 29 800
rect -29 -788 -17 788
rect 17 -788 29 788
rect -29 -800 29 -788
rect 229 788 287 800
rect 229 -788 241 788
rect 275 -788 287 788
rect 229 -800 287 -788
<< pdiffc >>
rect -275 -788 -241 788
rect -17 -788 17 788
rect 241 -788 275 788
<< poly >>
rect -229 800 -29 826
rect 29 800 229 826
rect -229 -826 -29 -800
rect 29 -826 229 -800
<< locali >>
rect -275 788 -241 804
rect -275 -804 -241 -788
rect -17 788 17 804
rect -17 -804 17 -788
rect 241 788 275 804
rect 241 -804 275 -788
<< viali >>
rect -275 -788 -241 788
rect -17 -788 17 788
rect 241 -788 275 788
<< metal1 >>
rect -281 788 -235 800
rect -281 -788 -275 788
rect -241 -788 -235 788
rect -281 -800 -235 -788
rect -23 788 23 800
rect -23 -788 -17 788
rect 17 -788 23 788
rect -23 -800 23 -788
rect 235 788 281 800
rect 235 -788 241 788
rect 275 -788 281 788
rect 235 -800 281 -788
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 8 l 1 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
