magic
tech sky130A
magscale 1 2
timestamp 1681046190
<< nwell >>
rect -387 -3262 387 3262
<< mvpmos >>
rect -129 -2964 -29 3036
rect 29 -2964 129 3036
<< mvpdiff >>
rect -187 3024 -129 3036
rect -187 -2952 -175 3024
rect -141 -2952 -129 3024
rect -187 -2964 -129 -2952
rect -29 3024 29 3036
rect -29 -2952 -17 3024
rect 17 -2952 29 3024
rect -29 -2964 29 -2952
rect 129 3024 187 3036
rect 129 -2952 141 3024
rect 175 -2952 187 3024
rect 129 -2964 187 -2952
<< mvpdiffc >>
rect -175 -2952 -141 3024
rect -17 -2952 17 3024
rect 141 -2952 175 3024
<< mvnsubdiff >>
rect -321 3184 321 3196
rect -321 3150 -213 3184
rect 213 3150 321 3184
rect -321 3138 321 3150
rect -321 3088 -263 3138
rect -321 -3088 -309 3088
rect -275 -3088 -263 3088
rect 263 3088 321 3138
rect -321 -3138 -263 -3088
rect 263 -3088 275 3088
rect 309 -3088 321 3088
rect 263 -3138 321 -3088
rect -321 -3150 321 -3138
rect -321 -3184 -213 -3150
rect 213 -3184 321 -3150
rect -321 -3196 321 -3184
<< mvnsubdiffcont >>
rect -213 3150 213 3184
rect -309 -3088 -275 3088
rect 275 -3088 309 3088
rect -213 -3184 213 -3150
<< poly >>
rect -129 3036 -29 3062
rect 29 3036 129 3062
rect -129 -3011 -29 -2964
rect -129 -3045 -113 -3011
rect -45 -3045 -29 -3011
rect -129 -3061 -29 -3045
rect 29 -3011 129 -2964
rect 29 -3045 45 -3011
rect 113 -3045 129 -3011
rect 29 -3061 129 -3045
<< polycont >>
rect -113 -3045 -45 -3011
rect 45 -3045 113 -3011
<< locali >>
rect -309 3150 -213 3184
rect 213 3150 309 3184
rect -309 3088 -275 3150
rect 275 3088 309 3150
rect -175 3024 -141 3040
rect -175 -2968 -141 -2952
rect -17 3024 17 3040
rect -17 -2968 17 -2952
rect 141 3024 175 3040
rect 141 -2968 175 -2952
rect -129 -3045 -113 -3011
rect -45 -3045 -29 -3011
rect 29 -3045 45 -3011
rect 113 -3045 129 -3011
rect -309 -3150 -275 -3088
rect 275 -3150 309 -3088
rect -309 -3184 -213 -3150
rect 213 -3184 309 -3150
<< viali >>
rect -175 -2952 -141 3024
rect -17 -2952 17 3024
rect 141 -2952 175 3024
rect -113 -3045 -45 -3011
rect 45 -3045 113 -3011
<< metal1 >>
rect -181 3024 -135 3036
rect -181 -2952 -175 3024
rect -141 -2952 -135 3024
rect -181 -2964 -135 -2952
rect -23 3024 23 3036
rect -23 -2952 -17 3024
rect 17 -2952 23 3024
rect -23 -2964 23 -2952
rect 135 3024 181 3036
rect 135 -2952 141 3024
rect 175 -2952 181 3024
rect 135 -2964 181 -2952
rect -125 -3011 -33 -3005
rect -125 -3045 -113 -3011
rect -45 -3045 -33 -3011
rect -125 -3051 -33 -3045
rect 33 -3011 125 -3005
rect 33 -3045 45 -3011
rect 113 -3045 125 -3011
rect 33 -3051 125 -3045
<< properties >>
string FIXED_BBOX -292 -3167 292 3167
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 30 l 0.50 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
