magic
tech sky130A
magscale 1 2
timestamp 1686989340
<< error_p >>
rect -194 -180 194 -114
rect -194 -283 -128 -180
rect -36 -283 36 -180
rect 128 -283 194 -180
rect -194 -349 194 -283
<< mvpdiff >>
rect -128 -237 -30 -180
rect -128 -271 -116 -237
rect -42 -271 -30 -237
rect -128 -283 -30 -271
rect 30 -237 128 -180
rect 30 -271 42 -237
rect 116 -271 128 -237
rect 30 -283 128 -271
<< mvpdiffc >>
rect -116 -271 -42 -237
rect 42 -271 116 -237
<< mvpdiffres >>
rect -128 186 128 284
rect -128 -180 -30 186
rect 30 -180 128 186
<< locali >>
rect -132 -271 -116 -237
rect -42 -271 -26 -237
rect 26 -271 42 -237
rect 116 -271 132 -237
<< properties >>
string gencell sky130_fd_pr__res_generic_pd__hv
string library sky130
string parameters w 0.488 l 2.1 m 1 nx 2 wmin 0.42 lmin 2.10 rho 197 val 2.217k dummy 0 dw 0.02 term 0.0 sterm 0.0 caplen 0.60 snake 1 guard 0 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
