magic
tech sky130A
magscale 1 2
timestamp 1686994090
<< nwell >>
rect 331 1860 4690 2280
rect 331 1833 4130 1860
rect 730 1820 4130 1833
rect 730 1200 3431 1820
rect 730 320 3440 1200
rect 4440 320 4690 1860
rect 730 140 4690 320
<< mvpmos >>
rect 2470 226 2550 250
<< mvpsubdiff >>
rect 1070 -1060 4200 -1010
rect 1070 -1260 1190 -1060
rect 4110 -1260 4200 -1060
rect 1070 -1310 4200 -1260
<< mvnsubdiff >>
rect 510 2140 4040 2200
rect 510 1960 610 2140
rect 1630 1960 1750 2140
rect 2760 1960 2920 2140
rect 3940 1960 4040 2140
rect 510 1900 4040 1960
<< mvpsubdiffcont >>
rect 1190 -1260 4110 -1060
<< mvnsubdiffcont >>
rect 610 1960 1630 2140
rect 1750 1960 2760 2140
rect 2920 1960 3940 2140
<< poly >>
rect 1840 1339 1897 1413
rect 1834 1329 1903 1339
rect 1834 1292 1850 1329
rect 1887 1292 1903 1329
rect 1834 1282 1903 1292
rect 2902 949 2959 1000
rect 3162 949 3219 1000
rect 2896 939 2965 949
rect 2896 902 2912 939
rect 2949 902 2965 939
rect 2896 892 2965 902
rect 3156 939 3225 949
rect 3156 902 3172 939
rect 3209 902 3225 939
rect 3156 892 3225 902
rect 1592 299 1649 350
rect 1842 299 1899 350
rect 1586 289 1655 299
rect 1586 242 1602 289
rect 1639 242 1655 289
rect 1586 232 1655 242
rect 1836 289 1905 299
rect 1836 242 1852 289
rect 1889 242 1905 289
rect 1836 232 1905 242
rect 952 149 1009 200
rect 1212 149 1269 200
rect 1696 178 1762 188
rect 1350 158 1416 168
rect 946 139 1015 149
rect 946 102 962 139
rect 999 102 1015 139
rect 946 92 1015 102
rect 1206 139 1275 149
rect 1206 102 1222 139
rect 1259 102 1275 139
rect 1350 124 1366 158
rect 1400 124 1416 158
rect 1696 144 1712 178
rect 1746 144 1762 178
rect 2222 149 2279 242
rect 2470 200 2550 226
rect 2812 219 2869 270
rect 3212 219 3269 270
rect 2806 209 2875 219
rect 2482 149 2539 200
rect 2806 162 2822 209
rect 2859 162 2875 209
rect 2806 152 2875 162
rect 3206 209 3275 219
rect 3206 162 3222 209
rect 3259 162 3275 209
rect 3206 152 3275 162
rect 3582 149 3639 200
rect 3842 149 3899 200
rect 4102 149 4159 200
rect 4352 149 4409 200
rect 1696 134 1762 144
rect 2216 139 2285 149
rect 1350 114 1416 124
rect 1206 92 1275 102
rect 1367 72 1399 114
rect 1713 92 1745 134
rect 2216 102 2232 139
rect 2269 102 2285 139
rect 2216 92 2285 102
rect 2476 139 2545 149
rect 2476 102 2492 139
rect 2529 102 2545 139
rect 2476 92 2545 102
rect 3576 139 3645 149
rect 3576 92 3592 139
rect 3629 92 3645 139
rect 1694 87 1773 92
rect 3576 82 3645 92
rect 3836 139 3905 149
rect 3836 92 3852 139
rect 3889 92 3905 139
rect 3836 82 3905 92
rect 4096 139 4165 149
rect 4096 92 4112 139
rect 4149 92 4165 139
rect 4096 82 4165 92
rect 4346 139 4415 149
rect 4346 92 4362 139
rect 4399 92 4415 139
rect 4346 82 4415 92
rect 1115 -2 1181 8
rect 1115 -36 1131 -2
rect 1165 -36 1181 -2
rect 1115 -46 1181 -36
rect 3576 -16 3642 -6
rect 1132 -88 1164 -46
rect 3576 -50 3592 -16
rect 3626 -50 3642 -16
rect 3576 -60 3642 -50
rect 3843 -16 3909 -6
rect 3843 -50 3859 -16
rect 3893 -50 3909 -16
rect 3843 -60 3909 -50
rect 4096 -16 4162 -6
rect 4096 -50 4112 -16
rect 4146 -50 4162 -16
rect 4096 -60 4162 -50
rect 4359 -16 4425 -6
rect 4359 -50 4375 -16
rect 4409 -50 4425 -16
rect 4359 -60 4425 -50
rect 3593 -102 3625 -60
rect 3860 -102 3892 -60
rect 4113 -102 4145 -60
rect 4376 -102 4408 -60
rect 3015 -242 3084 -232
rect 3015 -289 3031 -242
rect 3068 -289 3084 -242
rect 3015 -299 3084 -289
rect 3145 -242 3214 -232
rect 3145 -289 3161 -242
rect 3198 -289 3214 -242
rect 3145 -299 3214 -289
rect 3021 -350 3078 -299
rect 3151 -350 3208 -299
rect 2022 -842 2079 -791
rect 2016 -852 2085 -842
rect 2306 -844 2363 -793
rect 2672 -841 2729 -790
rect 1522 -903 1579 -860
rect 1712 -903 1769 -860
rect 2016 -899 2032 -852
rect 2069 -899 2085 -852
rect 1516 -913 1585 -903
rect 1516 -960 1532 -913
rect 1569 -960 1585 -913
rect 1516 -970 1585 -960
rect 1706 -913 1775 -903
rect 2016 -909 2085 -899
rect 2300 -854 2369 -844
rect 2300 -901 2316 -854
rect 2353 -901 2369 -854
rect 2300 -911 2369 -901
rect 2666 -851 2735 -841
rect 2666 -898 2682 -851
rect 2719 -898 2735 -851
rect 2666 -908 2735 -898
rect 1706 -960 1722 -913
rect 1759 -960 1775 -913
rect 1706 -970 1775 -960
<< polycont >>
rect 1850 1292 1887 1329
rect 2912 902 2949 939
rect 3172 902 3209 939
rect 1602 242 1639 289
rect 1852 242 1889 289
rect 962 102 999 139
rect 1222 102 1259 139
rect 1366 124 1400 158
rect 1712 144 1746 178
rect 2822 162 2859 209
rect 3222 162 3259 209
rect 2232 102 2269 139
rect 2492 102 2529 139
rect 3592 92 3629 139
rect 3852 92 3889 139
rect 4112 92 4149 139
rect 4362 92 4399 139
rect 1131 -36 1165 -2
rect 3592 -50 3626 -16
rect 3859 -50 3893 -16
rect 4112 -50 4146 -16
rect 4375 -50 4409 -16
rect 3031 -289 3068 -242
rect 3161 -289 3198 -242
rect 2032 -899 2069 -852
rect 1532 -960 1569 -913
rect 2316 -901 2353 -854
rect 2682 -898 2719 -851
rect 1722 -960 1759 -913
<< locali >>
rect 510 2140 4040 2200
rect 510 1960 610 2140
rect 1630 1960 1750 2140
rect 2760 1960 2920 2140
rect 3940 1960 4040 2140
rect 510 1900 4040 1960
rect 567 1096 639 1102
rect 567 1036 573 1096
rect 633 1036 639 1096
rect 1710 1095 1760 1495
rect 1850 1339 1887 1345
rect 1850 1276 1887 1282
rect 424 764 497 975
rect 567 824 639 1036
rect 2912 949 2949 955
rect 3172 949 3209 955
rect 2912 886 2949 892
rect 3172 886 3209 892
rect 671 764 715 766
rect 424 761 715 764
rect 424 721 671 761
rect 709 721 715 761
rect 424 716 715 721
rect 424 714 711 716
rect 424 596 497 714
rect 588 -820 660 662
rect 1602 299 1639 305
rect 1852 299 1889 305
rect 1602 226 1639 232
rect 1852 226 1889 232
rect 1712 178 1746 194
rect 1366 170 1400 174
rect 962 149 999 155
rect 1222 149 1259 155
rect 1405 144 1712 170
rect 1974 176 2008 379
rect 2930 290 3040 340
rect 2822 219 2859 225
rect 1746 144 1750 170
rect 1405 120 1750 144
rect 1788 142 2008 176
rect 2232 149 2269 155
rect 2492 149 2529 155
rect 1366 108 1400 120
rect 962 86 999 92
rect 1222 86 1259 92
rect 1131 -2 1165 14
rect 1788 7 1822 142
rect 2104 98 2138 109
rect 1907 64 2138 98
rect 2610 147 2680 150
rect 2610 113 2613 147
rect 2647 113 2680 147
rect 2822 146 2859 152
rect 2990 125 3040 290
rect 3222 219 3259 225
rect 3222 146 3259 152
rect 3592 149 3629 155
rect 3852 149 3889 155
rect 4112 149 4149 155
rect 4362 149 4399 155
rect 2610 110 2680 113
rect 2232 86 2269 92
rect 2492 86 2529 92
rect 2280 7 2360 10
rect 1989 -35 2070 5
rect 2280 -27 2283 7
rect 2317 -27 2360 7
rect 2280 -30 2360 -27
rect 1131 -52 1165 -36
rect 448 -906 477 -872
rect 2030 -570 2070 -35
rect 2030 -842 2070 -610
rect 2320 -710 2360 -30
rect 2640 -80 2680 110
rect 2935 75 3040 125
rect 3367 90 3582 140
rect 2935 -245 2985 75
rect 3367 -80 3407 90
rect 3639 90 3842 140
rect 3899 90 4102 140
rect 4159 90 4352 140
rect 4409 90 4410 140
rect 3592 76 3629 82
rect 3852 76 3889 82
rect 4112 76 4149 82
rect 4362 76 4399 82
rect 3592 -10 3626 0
rect 3859 -10 3893 0
rect 4112 -10 4146 0
rect 4375 -10 4409 0
rect 3630 -16 4409 -10
rect 3630 -50 3859 -16
rect 3893 -50 4112 -16
rect 4146 -50 4375 -16
rect 3592 -66 3626 -50
rect 3859 -66 3893 -50
rect 4112 -66 4146 -50
rect 4375 -66 4409 -50
rect 3080 -120 3407 -80
rect 3031 -232 3068 -226
rect 3161 -232 3198 -226
rect 2935 -295 3021 -245
rect 2935 -405 2985 -295
rect 3031 -305 3068 -299
rect 3161 -305 3198 -299
rect 2320 -838 2360 -750
rect 2316 -844 2360 -838
rect 2682 -841 2719 -835
rect 830 -920 880 -860
rect 1532 -903 1569 -897
rect 1722 -903 1759 -897
rect 1579 -962 1712 -912
rect 2032 -915 2069 -909
rect 2316 -917 2353 -911
rect 2682 -914 2719 -908
rect 1532 -976 1569 -970
rect 1722 -976 1759 -970
rect 1070 -1060 4200 -1010
rect 1070 -1260 1190 -1060
rect 4110 -1260 4200 -1060
rect 1070 -1310 4200 -1260
<< viali >>
rect 610 1960 1630 2140
rect 1750 1960 2760 2140
rect 2920 1960 3940 2140
rect 573 1036 633 1096
rect 1840 1329 1897 1339
rect 1840 1292 1850 1329
rect 1850 1292 1887 1329
rect 1887 1292 1897 1329
rect 1840 1282 1897 1292
rect 2902 939 2959 949
rect 2902 902 2912 939
rect 2912 902 2949 939
rect 2949 902 2959 939
rect 2902 892 2959 902
rect 3162 939 3219 949
rect 3162 902 3172 939
rect 3172 902 3209 939
rect 3209 902 3219 939
rect 3162 892 3219 902
rect 671 721 709 761
rect 1592 289 1649 299
rect 1592 242 1602 289
rect 1602 242 1639 289
rect 1639 242 1649 289
rect 1592 232 1649 242
rect 1842 289 1899 299
rect 1842 242 1852 289
rect 1852 242 1889 289
rect 1889 242 1899 289
rect 1842 232 1899 242
rect 1355 158 1405 170
rect 952 139 1009 149
rect 952 102 962 139
rect 962 102 999 139
rect 999 102 1009 139
rect 952 92 1009 102
rect 1212 139 1269 149
rect 1212 102 1222 139
rect 1222 102 1259 139
rect 1259 102 1269 139
rect 1355 124 1366 158
rect 1366 124 1400 158
rect 1400 124 1405 158
rect 1712 144 1746 178
rect 1355 120 1405 124
rect 2812 209 2869 219
rect 2812 162 2822 209
rect 2822 162 2859 209
rect 2859 162 2869 209
rect 2812 152 2869 162
rect 1212 92 1269 102
rect 2104 109 2138 143
rect 1873 64 1907 98
rect 2222 139 2279 149
rect 2222 102 2232 139
rect 2232 102 2269 139
rect 2269 102 2279 139
rect 2222 92 2279 102
rect 2482 139 2539 149
rect 2482 102 2492 139
rect 2492 102 2529 139
rect 2529 102 2539 139
rect 2613 113 2647 147
rect 3212 209 3269 219
rect 3212 162 3222 209
rect 3222 162 3259 209
rect 3259 162 3269 209
rect 3212 152 3269 162
rect 2482 92 2539 102
rect 1131 -36 1165 -2
rect 1949 -35 1989 5
rect 2283 -27 2317 7
rect 414 -906 448 -872
rect 588 -892 660 -820
rect 2030 -610 2070 -570
rect 2640 -120 2680 -80
rect 3582 139 3639 149
rect 3582 92 3592 139
rect 3592 92 3629 139
rect 3629 92 3639 139
rect 3582 82 3639 92
rect 3842 139 3899 149
rect 3842 92 3852 139
rect 3852 92 3889 139
rect 3889 92 3899 139
rect 3842 82 3899 92
rect 4102 139 4159 149
rect 4102 92 4112 139
rect 4112 92 4149 139
rect 4149 92 4159 139
rect 4102 82 4159 92
rect 4352 139 4409 149
rect 4352 92 4362 139
rect 4362 92 4399 139
rect 4399 92 4409 139
rect 4352 82 4409 92
rect 3590 -16 3630 -10
rect 3590 -50 3592 -16
rect 3592 -50 3626 -16
rect 3626 -50 3630 -16
rect 3859 -50 3893 -16
rect 4112 -50 4146 -16
rect 4375 -50 4409 -16
rect 3046 -120 3080 -80
rect 3021 -242 3078 -232
rect 3021 -289 3031 -242
rect 3031 -289 3068 -242
rect 3068 -289 3078 -242
rect 3021 -299 3078 -289
rect 3151 -242 3208 -232
rect 3151 -289 3161 -242
rect 3161 -289 3198 -242
rect 3198 -289 3208 -242
rect 3151 -299 3208 -289
rect 2320 -750 2360 -710
rect 2022 -852 2079 -842
rect 880 -920 940 -860
rect 2022 -899 2032 -852
rect 2032 -899 2069 -852
rect 2069 -899 2079 -852
rect 1522 -913 1579 -903
rect 1522 -960 1532 -913
rect 1532 -960 1569 -913
rect 1569 -960 1579 -913
rect 1522 -970 1579 -960
rect 1712 -913 1769 -903
rect 2022 -909 2079 -899
rect 2306 -854 2363 -844
rect 2306 -901 2316 -854
rect 2316 -901 2353 -854
rect 2353 -901 2363 -854
rect 1712 -960 1722 -913
rect 1722 -960 1759 -913
rect 1759 -960 1769 -913
rect 2306 -911 2363 -901
rect 2672 -851 2729 -841
rect 2672 -898 2682 -851
rect 2682 -898 2719 -851
rect 2719 -898 2729 -851
rect 2672 -908 2729 -898
rect 1712 -970 1769 -960
rect 1190 -1260 4110 -1060
<< metal1 >>
rect 510 2140 4560 2200
rect 510 1960 610 2140
rect 1630 1960 1750 2140
rect 2760 1960 2920 2140
rect 3940 1960 4560 2140
rect 510 1900 4560 1960
rect 567 1096 639 1900
rect 1070 1800 1120 1900
rect 1330 1596 1370 1860
rect 1970 1790 2020 1900
rect 2350 1800 2400 1900
rect 3030 1780 3080 1900
rect 3460 1790 3510 1900
rect 3970 1800 4020 1900
rect 4490 1800 4540 1900
rect 1318 1544 1324 1596
rect 1376 1590 1382 1596
rect 1376 1550 1383 1590
rect 1376 1544 1382 1550
rect 1834 1339 1903 1351
rect 1506 1282 1512 1339
rect 1569 1282 1840 1339
rect 1900 1282 1906 1339
rect 1834 1270 1903 1282
rect 567 1036 573 1096
rect 633 1036 639 1096
rect 567 1024 639 1036
rect 2770 835 2820 1040
rect 2896 958 2965 961
rect 2888 952 2965 958
rect 2945 949 2976 952
rect 2959 937 2976 949
rect 3156 949 3225 961
rect 3156 937 3162 949
rect 2959 904 3162 937
rect 2959 895 2976 904
rect 2888 892 2902 895
rect 2959 892 2965 895
rect 2888 889 2965 892
rect 2896 880 2965 889
rect 3156 892 3162 904
rect 3219 937 3225 949
rect 3219 904 3230 937
rect 3219 892 3225 904
rect 3156 880 3225 892
rect 3290 845 3340 1135
rect 2735 785 2820 835
rect 3145 795 3340 845
rect 665 767 717 773
rect 659 715 665 767
rect 717 715 721 767
rect 665 709 717 715
rect 2735 412 2785 785
rect 3145 626 3195 795
rect 3138 574 3144 626
rect 3196 574 3202 626
rect 2734 406 2786 412
rect 1206 272 1212 329
rect 1269 272 1275 329
rect 1457 290 1497 400
rect 2734 348 2786 354
rect 1586 299 1655 311
rect 824 137 857 256
rect 1212 161 1269 272
rect 1457 250 1510 290
rect 1586 287 1592 299
rect 1349 176 1411 182
rect 946 149 1015 161
rect 946 137 952 149
rect 824 104 952 137
rect 824 -733 857 104
rect 946 92 952 104
rect 1009 137 1015 149
rect 1206 149 1275 161
rect 1206 137 1212 149
rect 1009 104 1212 137
rect 1009 92 1015 104
rect 946 80 1015 92
rect 1206 92 1212 104
rect 1269 92 1275 149
rect 1343 124 1349 176
rect 1411 171 1417 176
rect 1411 124 1420 171
rect 1343 120 1355 124
rect 1405 120 1420 124
rect 1343 114 1420 120
rect 1351 113 1420 114
rect 1360 112 1406 113
rect 1206 80 1275 92
rect 1088 0 1094 12
rect 1030 -40 1094 0
rect 1146 11 1152 12
rect 1146 -2 1185 11
rect 1165 -36 1185 -2
rect 1299 -31 1305 21
rect 1357 -31 1363 21
rect 1470 0 1510 250
rect 1580 244 1592 287
rect 1649 287 1655 299
rect 1836 299 1905 311
rect 1836 287 1842 299
rect 1649 244 1660 287
rect 1830 244 1842 287
rect 1586 232 1592 244
rect 1649 232 1655 244
rect 1586 220 1655 232
rect 1836 232 1842 244
rect 1899 287 1905 299
rect 1899 244 1910 287
rect 1899 232 1905 244
rect 1836 220 1905 232
rect 1697 178 1766 191
rect 1697 144 1712 178
rect 1746 144 1766 178
rect 1850 190 1890 220
rect 1850 150 2070 190
rect 2104 155 2137 256
rect 1697 133 1766 144
rect 1706 132 1752 133
rect 1867 107 1913 110
rect 1858 55 1864 107
rect 1916 55 1922 107
rect 1867 52 1913 55
rect 1943 11 1995 17
rect 1146 -40 1185 -36
rect 1030 -150 1070 -40
rect 1116 -47 1185 -40
rect 1125 -48 1171 -47
rect 1314 -92 1348 -31
rect 1937 -41 1943 11
rect 1995 -41 2001 11
rect 2030 10 2070 150
rect 2098 143 2144 155
rect 2098 109 2104 143
rect 2138 137 2144 143
rect 2216 149 2285 161
rect 2216 137 2222 149
rect 2138 109 2222 137
rect 2098 104 2222 109
rect 2098 97 2144 104
rect 2216 92 2222 104
rect 2279 137 2285 149
rect 2476 149 2545 161
rect 2610 159 2650 240
rect 2806 222 2875 231
rect 2806 219 2876 222
rect 2806 207 2812 219
rect 2869 216 2876 219
rect 2800 164 2812 207
rect 3206 219 3275 231
rect 3206 210 3212 219
rect 2876 164 3212 210
rect 2476 137 2482 149
rect 2279 104 2482 137
rect 2279 92 2285 104
rect 2216 80 2285 92
rect 2476 92 2482 104
rect 2539 92 2545 149
rect 2607 147 2653 159
rect 2607 113 2613 147
rect 2647 113 2653 147
rect 2806 152 2812 164
rect 2869 160 3212 164
rect 2869 158 2876 160
rect 2869 152 2875 158
rect 2806 140 2875 152
rect 3206 152 3212 160
rect 3269 207 3275 219
rect 3269 164 3280 207
rect 3269 152 3275 164
rect 3206 140 3275 152
rect 2607 101 2653 113
rect 2476 80 2545 92
rect 3310 70 3350 310
rect 3576 149 3645 161
rect 3576 137 3582 149
rect 3570 94 3582 137
rect 3576 82 3582 94
rect 3639 137 3645 149
rect 3639 94 3650 137
rect 3720 136 3770 250
rect 3836 149 3905 161
rect 3836 137 3842 149
rect 3639 82 3645 94
rect 3713 84 3719 136
rect 3771 84 3777 136
rect 3830 94 3842 137
rect 3576 70 3645 82
rect 3260 30 3350 70
rect 2277 10 2323 19
rect 2030 7 2323 10
rect 2030 -27 2283 7
rect 2317 -27 2323 7
rect 2030 -30 2323 -27
rect 1943 -47 1995 -41
rect 2030 -51 2070 -30
rect 2277 -39 2323 -30
rect 3260 -10 3300 30
rect 3584 -3 3636 2
rect 3577 -10 3646 -3
rect 3260 -50 3590 -10
rect 3630 -50 3646 -10
rect 2194 -74 2246 -68
rect 1630 -134 1670 -80
rect 2434 -74 2486 -68
rect 2634 -74 2686 -68
rect 3034 -74 3086 -68
rect 2246 -120 2434 -80
rect 2194 -132 2246 -126
rect 2628 -126 2634 -74
rect 2686 -126 2692 -74
rect 3086 -126 3092 -74
rect 2434 -132 2486 -126
rect 2634 -132 2686 -126
rect 3034 -132 3086 -126
rect 1618 -140 1624 -134
rect 1616 -180 1624 -140
rect 1618 -186 1624 -180
rect 1676 -186 1682 -134
rect 2304 -184 2356 -178
rect 1630 -240 1670 -186
rect 1905 -235 2304 -185
rect 1460 -460 1510 -340
rect 1782 -456 1830 -300
rect 1905 -425 1955 -235
rect 2304 -242 2356 -236
rect 3015 -232 3084 -220
rect 3015 -244 3021 -232
rect 2160 -325 2585 -275
rect 3010 -287 3021 -244
rect 3015 -299 3021 -287
rect 3078 -240 3084 -232
rect 3145 -232 3214 -220
rect 3145 -240 3151 -232
rect 3078 -290 3151 -240
rect 3078 -299 3084 -290
rect 3015 -311 3084 -299
rect 3145 -299 3151 -290
rect 3208 -244 3214 -232
rect 3208 -287 3220 -244
rect 3208 -299 3214 -287
rect 3145 -311 3214 -299
rect 2160 -380 2210 -325
rect 2418 -466 2424 -414
rect 2476 -466 2482 -414
rect 3260 -430 3300 -50
rect 3577 -61 3646 -50
rect 3584 -62 3636 -61
rect 3720 -150 3770 84
rect 3836 82 3842 94
rect 3899 137 3905 149
rect 4096 149 4165 161
rect 4096 137 4102 149
rect 3899 94 3910 137
rect 4090 94 4102 137
rect 3899 82 3905 94
rect 3836 70 3905 82
rect 4096 82 4102 94
rect 4159 137 4165 149
rect 4159 94 4170 137
rect 4235 136 4285 265
rect 4346 149 4415 161
rect 4346 137 4352 149
rect 4159 82 4165 94
rect 4228 84 4234 136
rect 4286 84 4292 136
rect 4340 94 4352 137
rect 4096 70 4165 82
rect 3844 -16 3913 -3
rect 3844 -50 3859 -16
rect 3893 -50 3913 -16
rect 3844 -61 3913 -50
rect 4097 -16 4166 -3
rect 4097 -50 4112 -16
rect 4146 -50 4166 -16
rect 4097 -61 4166 -50
rect 3853 -62 3899 -61
rect 4106 -62 4152 -61
rect 4240 -150 4290 84
rect 4346 82 4352 94
rect 4409 137 4415 149
rect 4409 94 4420 137
rect 4409 82 4415 94
rect 4346 70 4415 82
rect 4360 -16 4429 -3
rect 4360 -50 4375 -16
rect 4409 -50 4429 -16
rect 4360 -61 4429 -50
rect 4369 -62 4415 -61
rect 2024 -564 2076 -558
rect 2018 -616 2024 -564
rect 2076 -616 2082 -564
rect 2425 -575 2475 -466
rect 3730 -564 3770 -150
rect 3718 -616 3724 -564
rect 3776 -616 3782 -564
rect 2024 -622 2076 -616
rect 2314 -704 2366 -698
rect 414 -766 857 -733
rect 2308 -756 2314 -704
rect 2366 -756 2372 -704
rect 2314 -762 2366 -756
rect 414 -866 447 -766
rect 576 -820 672 -814
rect 402 -872 460 -866
rect 402 -906 414 -872
rect 448 -906 460 -872
rect 576 -892 588 -820
rect 660 -892 672 -820
rect 576 -898 672 -892
rect 874 -860 946 -848
rect 402 -912 460 -906
rect 588 -1043 660 -898
rect 874 -920 880 -860
rect 940 -920 946 -860
rect 874 -932 946 -920
rect 880 -1043 940 -932
rect 1190 -1010 1230 -890
rect 1314 -904 1366 -898
rect 1516 -903 1585 -891
rect 1516 -910 1522 -903
rect 1366 -950 1522 -910
rect 1314 -962 1366 -956
rect 1510 -958 1522 -950
rect 1516 -970 1522 -958
rect 1579 -915 1585 -903
rect 1579 -958 1590 -915
rect 1579 -970 1585 -958
rect 1516 -982 1585 -970
rect 1630 -1010 1670 -780
rect 2016 -842 2085 -830
rect 2016 -854 2022 -842
rect 1706 -903 1775 -891
rect 2010 -897 2022 -854
rect 1706 -915 1712 -903
rect 1700 -958 1712 -915
rect 1706 -970 1712 -958
rect 1769 -907 1775 -903
rect 1925 -903 1977 -897
rect 1769 -950 1925 -907
rect 1769 -958 1780 -950
rect 2016 -909 2022 -897
rect 2079 -854 2085 -842
rect 2300 -844 2369 -832
rect 2079 -897 2090 -854
rect 2300 -856 2306 -844
rect 2079 -909 2085 -897
rect 2294 -899 2306 -856
rect 2016 -921 2085 -909
rect 2300 -911 2306 -899
rect 2363 -856 2369 -844
rect 2666 -841 2735 -829
rect 2363 -899 2374 -856
rect 2363 -911 2369 -899
rect 2509 -900 2515 -848
rect 2567 -853 2573 -848
rect 2666 -853 2672 -841
rect 2567 -896 2672 -853
rect 2567 -900 2573 -896
rect 2300 -923 2369 -911
rect 2666 -908 2672 -896
rect 2729 -853 2735 -841
rect 2729 -896 2740 -853
rect 2729 -908 2735 -896
rect 2666 -920 2735 -908
rect 1769 -970 1775 -958
rect 1925 -961 1977 -955
rect 1706 -982 1775 -970
rect 2800 -1010 2850 -715
rect 3090 -1010 3140 -760
rect 3460 -1010 3510 -826
rect 3980 -1010 4030 -816
rect 1070 -1043 4200 -1010
rect 588 -1055 4200 -1043
rect 4490 -1055 4540 -786
rect 588 -1060 4540 -1055
rect 588 -1115 1190 -1060
rect 1070 -1260 1190 -1115
rect 4110 -1105 4540 -1060
rect 4110 -1260 4200 -1105
rect 1070 -1310 4200 -1260
<< via1 >>
rect 610 1960 1630 2140
rect 1750 1960 2760 2140
rect 2920 1960 3940 2140
rect 1324 1544 1376 1596
rect 1512 1282 1569 1339
rect 1843 1282 1897 1339
rect 1897 1282 1900 1339
rect 2888 949 2945 952
rect 2888 895 2902 949
rect 2902 895 2945 949
rect 665 761 717 767
rect 665 721 671 761
rect 671 721 709 761
rect 709 721 717 761
rect 665 715 717 721
rect 3144 574 3196 626
rect 1212 272 1269 329
rect 2734 354 2786 406
rect 1349 170 1411 176
rect 1349 124 1355 170
rect 1355 124 1405 170
rect 1405 124 1411 170
rect 1094 -2 1146 12
rect 1094 -36 1131 -2
rect 1131 -36 1146 -2
rect 1305 -31 1357 21
rect 1594 244 1646 296
rect 1864 98 1916 107
rect 1864 64 1873 98
rect 1873 64 1907 98
rect 1907 64 1916 98
rect 1864 55 1916 64
rect 1094 -40 1146 -36
rect 1943 5 1995 11
rect 1943 -35 1949 5
rect 1949 -35 1989 5
rect 1989 -35 1995 5
rect 1943 -41 1995 -35
rect 2824 164 2869 216
rect 2869 164 2876 216
rect 3719 84 3771 136
rect 2194 -126 2246 -74
rect 2434 -126 2486 -74
rect 2634 -80 2686 -74
rect 2634 -120 2640 -80
rect 2640 -120 2680 -80
rect 2680 -120 2686 -80
rect 2634 -126 2686 -120
rect 3034 -80 3086 -74
rect 3034 -120 3046 -80
rect 3046 -120 3080 -80
rect 3080 -120 3086 -80
rect 3034 -126 3086 -120
rect 1624 -186 1676 -134
rect 2304 -236 2356 -184
rect 2424 -466 2476 -414
rect 4234 84 4286 136
rect 2024 -570 2076 -564
rect 2024 -610 2030 -570
rect 2030 -610 2070 -570
rect 2070 -610 2076 -570
rect 2024 -616 2076 -610
rect 3724 -616 3776 -564
rect 2314 -710 2366 -704
rect 2314 -750 2320 -710
rect 2320 -750 2360 -710
rect 2360 -750 2366 -710
rect 2314 -756 2366 -750
rect 1314 -956 1366 -904
rect 1925 -955 1977 -903
rect 2515 -900 2567 -848
rect 1190 -1260 4110 -1060
<< metal2 >>
rect 510 2140 4040 2200
rect 510 1960 610 2140
rect 1630 1960 1750 2140
rect 2760 1960 2920 2140
rect 3940 1960 4040 2140
rect 510 1900 4040 1960
rect 923 1652 3081 1702
rect 659 715 665 767
rect 717 766 723 767
rect 923 766 973 1652
rect 1324 1596 1376 1602
rect 717 716 973 766
rect 1100 1550 1324 1590
rect 717 715 723 716
rect 1100 18 1140 1550
rect 1324 1538 1376 1544
rect 1512 1339 1569 1345
rect 1212 1282 1512 1339
rect 1212 329 1269 1282
rect 1512 1276 1569 1282
rect 1843 1339 1900 1345
rect 1900 1282 2945 1339
rect 1843 1276 1900 1282
rect 2888 952 2945 1282
rect 2882 895 2888 952
rect 2945 895 2951 952
rect 3031 782 3081 1652
rect 2825 732 3081 782
rect 2825 585 2875 732
rect 1212 266 1269 272
rect 1355 535 2875 585
rect 3144 626 3196 632
rect 3144 568 3196 574
rect 1355 176 1405 535
rect 2728 354 2734 406
rect 2786 354 2792 406
rect 1588 244 1594 296
rect 1646 290 1652 296
rect 1646 250 1988 290
rect 1646 244 1652 250
rect 1343 124 1349 176
rect 1411 124 1417 176
rect 1864 110 1916 113
rect 1860 107 1920 110
rect 1860 88 1864 107
rect 1314 55 1864 88
rect 1916 55 1920 107
rect 1314 54 1920 55
rect 1314 27 1360 54
rect 1860 50 1920 54
rect 1864 49 1916 50
rect 1305 21 1360 27
rect 1094 12 1146 18
rect 1146 -40 1260 0
rect 1357 10 1360 21
rect 1948 11 1988 250
rect 2735 35 2785 354
rect 2825 216 2875 535
rect 2818 164 2824 216
rect 2876 164 2882 216
rect 1305 -37 1357 -31
rect 1094 -46 1146 -40
rect 1220 -500 1260 -40
rect 1937 -41 1943 11
rect 1995 -41 2001 11
rect 2305 -15 2785 35
rect 2188 -80 2194 -74
rect 1880 -120 2194 -80
rect 1624 -134 1676 -128
rect 1880 -140 1920 -120
rect 2188 -126 2194 -120
rect 2246 -126 2252 -74
rect 1676 -180 1920 -140
rect 2305 -184 2355 -15
rect 2634 -74 2686 -68
rect 2428 -126 2434 -74
rect 2486 -80 2492 -74
rect 2486 -120 2634 -80
rect 2486 -126 2492 -120
rect 3028 -80 3034 -74
rect 2686 -120 3034 -80
rect 3028 -126 3034 -120
rect 3086 -126 3092 -74
rect 2634 -132 2686 -126
rect 1624 -192 1676 -186
rect 2298 -236 2304 -184
rect 2356 -236 2362 -184
rect 3145 -247 3195 568
rect 3719 136 3771 142
rect 4234 136 4286 142
rect 3771 85 4234 135
rect 3719 78 3771 84
rect 4286 85 4541 135
rect 4234 78 4286 84
rect 4491 49 4541 85
rect 4491 -1 4689 49
rect 2425 -297 3195 -247
rect 2425 -408 2475 -297
rect 2424 -414 2476 -408
rect 2424 -472 2476 -466
rect 1220 -540 1360 -500
rect 1320 -904 1360 -540
rect 2024 -564 2076 -558
rect 3724 -564 3776 -558
rect 2076 -610 3724 -570
rect 2024 -622 2076 -616
rect 3724 -622 3776 -616
rect 2314 -704 2366 -698
rect 2366 -750 4696 -710
rect 2314 -762 2366 -756
rect 2515 -848 2567 -842
rect 2189 -895 2515 -852
rect 1308 -956 1314 -904
rect 1366 -956 1372 -904
rect 1919 -955 1925 -903
rect 1977 -908 1983 -903
rect 2189 -908 2232 -895
rect 2515 -906 2567 -900
rect 1977 -951 2232 -908
rect 1977 -955 1983 -951
rect 1070 -1060 4200 -1010
rect 1070 -1260 1190 -1060
rect 4110 -1260 4200 -1060
rect 1070 -1310 4200 -1260
<< via2 >>
rect 610 1960 1630 2140
rect 1750 1960 2760 2140
rect 2920 1960 3940 2140
rect 1190 -1260 4110 -1060
<< metal3 >>
rect 272 2140 4741 2200
rect 272 1960 610 2140
rect 1630 1960 1750 2140
rect 2760 1960 2920 2140
rect 3940 1960 4741 2140
rect 272 1900 4741 1960
rect 272 -1060 4741 -1010
rect 272 -1260 1190 -1060
rect 4110 -1260 4741 -1060
rect 272 -1310 4741 -1260
use sky130_fd_pr__nfet_g5v0d10v5_4DV7XU  sky130_fd_pr__nfet_g5v0d10v5_4DV7XU_0
timestamp 1686988006
transform 1 0 4001 0 1 -528
box -545 -426 545 426
use sky130_fd_pr__nfet_g5v0d10v5_GEEYVT  sky130_fd_pr__nfet_g5v0d10v5_GEEYVT_0
timestamp 1686986091
transform 1 0 2187 0 1 -574
box -287 -226 287 226
use sky130_fd_pr__nfet_g5v0d10v5_N5C7ZL  sky130_fd_pr__nfet_g5v0d10v5_N5C7ZL_0
timestamp 1686986091
transform 1 0 1647 0 1 -634
box -187 -226 187 226
use sky130_fd_pr__nfet_g5v0d10v5_N5C7ZL  sky130_fd_pr__nfet_g5v0d10v5_N5C7ZL_1
timestamp 1686986091
transform 1 0 3117 0 1 -574
box -187 -226 187 226
use sky130_fd_pr__nfet_g5v0d10v5_NY97Z6  sky130_fd_pr__nfet_g5v0d10v5_NY97Z6_0
timestamp 1686986091
transform 1 0 1726 0 1 -134
box -108 -226 108 226
use sky130_fd_pr__nfet_g5v0d10v5_NY97Z6  sky130_fd_pr__nfet_g5v0d10v5_NY97Z6_1
timestamp 1686986091
transform 1 0 1408 0 1 -154
box -108 -226 108 226
use sky130_fd_pr__nfet_g5v0d10v5_TNBBPH  sky130_fd_pr__nfet_g5v0d10v5_TNBBPH_0
timestamp 1686986870
transform 1 0 1130 0 1 -514
box -108 -426 108 426
use sky130_fd_pr__nfet_g5v0d10v5_UEV7X2  sky130_fd_pr__nfet_g5v0d10v5_UEV7X2_0
timestamp 1686986091
transform 1 0 2698 0 1 -364
box -158 -426 158 426
use sky130_fd_pr__pfet_g5v0d10v5_5HRSW2  sky130_fd_pr__pfet_g5v0d10v5_5HRSW2_0
timestamp 1686986091
transform 1 0 1864 0 1 1616
box -224 -266 224 266
use sky130_fd_pr__pfet_g5v0d10v5_BHVYLS  sky130_fd_pr__pfet_g5v0d10v5_BHVYLS_0
timestamp 1686986091
transform 1 0 3053 0 1 1426
box -353 -466 353 466
use sky130_fd_pr__pfet_g5v0d10v5_BHVYLS  sky130_fd_pr__pfet_g5v0d10v5_BHVYLS_1
timestamp 1686986091
transform 1 0 1733 0 1 776
box -353 -466 353 466
use sky130_fd_pr__pfet_g5v0d10v5_EH58LG  sky130_fd_pr__pfet_g5v0d10v5_EH58LG_0
timestamp 1686986091
transform 1 0 4001 0 1 1024
box -611 -866 611 866
use sky130_fd_pr__pfet_g5v0d10v5_EHVYLG  sky130_fd_pr__pfet_g5v0d10v5_EHVYLG_0
timestamp 1686986091
transform 1 0 1093 0 1 1026
box -353 -866 353 866
use sky130_fd_pr__pfet_g5v0d10v5_EHVYLG  sky130_fd_pr__pfet_g5v0d10v5_EHVYLG_1
timestamp 1686986091
transform 1 0 2373 0 1 1026
box -353 -866 353 866
use sky130_fd_pr__pfet_g5v0d10v5_SVVZZ7  sky130_fd_pr__pfet_g5v0d10v5_SVVZZ7_0
timestamp 1686986091
transform 1 0 3254 0 1 492
box -174 -266 174 266
use sky130_fd_pr__pfet_g5v0d10v5_SVVZZ7  sky130_fd_pr__pfet_g5v0d10v5_SVVZZ7_1
timestamp 1686986091
transform 1 0 2844 0 1 492
box -174 -266 174 266
use sky130_fd_pr__res_generic_nd__hv_CGSFZ8  sky130_fd_pr__res_generic_nd__hv_CGSFZ8_0
timestamp 1686990252
transform -1 0 535 0 -1 372
box -130 -283 130 284
use sky130_fd_pr__res_generic_nd__hv_FHMM3Y  sky130_fd_pr__res_generic_nd__hv_FHMM3Y_0
timestamp 1686993383
transform 1 0 530 0 1 1293
box -118 -473 118 474
use sky130_fd_pr__res_generic_nd__hv_FMMP3Y  sky130_fd_pr__res_generic_nd__hv_FMMP3Y_0
timestamp 1686987678
transform 1 0 652 0 1 -447
box -262 -473 262 474
<< labels >>
flabel metal3 s 340 -1190 340 -1190 0 FreeSans 640 0 0 0 VSSA
flabel metal2 s 4668 -732 4668 -732 0 FreeSans 800 0 0 0 VIN
flabel metal2 s 4660 26 4660 26 0 FreeSans 800 0 0 0 VOUT
flabel metal3 s 391 2063 391 2063 0 FreeSans 640 0 0 0 VDDA
<< end >>
