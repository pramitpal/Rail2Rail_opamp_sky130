magic
tech sky130A
timestamp 1678605198
<< nmos >>
rect -10 -400 10 400
<< ndiff >>
rect -39 394 -10 400
rect -39 -394 -33 394
rect -16 -394 -10 394
rect -39 -400 -10 -394
rect 10 394 39 400
rect 10 -394 16 394
rect 33 -394 39 394
rect 10 -400 39 -394
<< ndiffc >>
rect -33 -394 -16 394
rect 16 -394 33 394
<< poly >>
rect -10 400 10 413
rect -10 -413 10 -400
<< locali >>
rect -33 394 -16 402
rect -33 -402 -16 -394
rect 16 394 33 402
rect 16 -402 33 -394
<< viali >>
rect -33 -394 -16 394
rect 16 -394 33 394
<< metal1 >>
rect -36 394 -13 400
rect -36 -394 -33 394
rect -16 -394 -13 394
rect -36 -400 -13 -394
rect 13 394 36 400
rect 13 -394 16 394
rect 33 -394 36 394
rect 13 -400 36 -394
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 8 l 0.2 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
