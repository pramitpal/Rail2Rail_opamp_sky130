magic
tech sky130A
magscale 1 2
timestamp 1681052864
<< error_p >>
rect -411 1098 411 1102
rect -411 -1030 -381 1098
rect -345 1032 345 1036
rect -345 -964 -315 1032
rect 315 -964 345 1032
rect 381 -1030 411 1098
<< nwell >>
rect -381 -1064 381 1098
<< mvpmos >>
rect -287 -964 -187 1036
rect -129 -964 -29 1036
rect 29 -964 129 1036
rect 187 -964 287 1036
<< mvpdiff >>
rect -345 1024 -287 1036
rect -345 -952 -333 1024
rect -299 -952 -287 1024
rect -345 -964 -287 -952
rect -187 1024 -129 1036
rect -187 -952 -175 1024
rect -141 -952 -129 1024
rect -187 -964 -129 -952
rect -29 1024 29 1036
rect -29 -952 -17 1024
rect 17 -952 29 1024
rect -29 -964 29 -952
rect 129 1024 187 1036
rect 129 -952 141 1024
rect 175 -952 187 1024
rect 129 -964 187 -952
rect 287 1024 345 1036
rect 287 -952 299 1024
rect 333 -952 345 1024
rect 287 -964 345 -952
<< mvpdiffc >>
rect -333 -952 -299 1024
rect -175 -952 -141 1024
rect -17 -952 17 1024
rect 141 -952 175 1024
rect 299 -952 333 1024
<< poly >>
rect -287 1036 -187 1062
rect -129 1036 -29 1062
rect 29 1036 129 1062
rect 187 1036 287 1062
rect -287 -1011 -187 -964
rect -287 -1045 -271 -1011
rect -203 -1045 -187 -1011
rect -287 -1061 -187 -1045
rect -129 -1011 -29 -964
rect -129 -1045 -113 -1011
rect -45 -1045 -29 -1011
rect -129 -1061 -29 -1045
rect 29 -1011 129 -964
rect 29 -1045 45 -1011
rect 113 -1045 129 -1011
rect 29 -1061 129 -1045
rect 187 -1011 287 -964
rect 187 -1045 203 -1011
rect 271 -1045 287 -1011
rect 187 -1061 287 -1045
<< polycont >>
rect -271 -1045 -203 -1011
rect -113 -1045 -45 -1011
rect 45 -1045 113 -1011
rect 203 -1045 271 -1011
<< locali >>
rect -333 1024 -299 1040
rect -333 -968 -299 -952
rect -175 1024 -141 1040
rect -175 -968 -141 -952
rect -17 1024 17 1040
rect -17 -968 17 -952
rect 141 1024 175 1040
rect 141 -968 175 -952
rect 299 1024 333 1040
rect 299 -968 333 -952
rect -287 -1045 -271 -1011
rect -203 -1045 -187 -1011
rect -129 -1045 -113 -1011
rect -45 -1045 -29 -1011
rect 29 -1045 45 -1011
rect 113 -1045 129 -1011
rect 187 -1045 203 -1011
rect 271 -1045 287 -1011
<< viali >>
rect -333 -952 -299 1024
rect -175 -952 -141 1024
rect -17 -952 17 1024
rect 141 -952 175 1024
rect 299 -952 333 1024
rect -271 -1045 -203 -1011
rect -113 -1045 -45 -1011
rect 45 -1045 113 -1011
rect 203 -1045 271 -1011
<< metal1 >>
rect -339 1024 -293 1036
rect -339 -952 -333 1024
rect -299 -952 -293 1024
rect -339 -964 -293 -952
rect -181 1024 -135 1036
rect -181 -952 -175 1024
rect -141 -952 -135 1024
rect -181 -964 -135 -952
rect -23 1024 23 1036
rect -23 -952 -17 1024
rect 17 -952 23 1024
rect -23 -964 23 -952
rect 135 1024 181 1036
rect 135 -952 141 1024
rect 175 -952 181 1024
rect 135 -964 181 -952
rect 293 1024 339 1036
rect 293 -952 299 1024
rect 333 -952 339 1024
rect 293 -964 339 -952
rect -283 -1011 -191 -1005
rect -283 -1045 -271 -1011
rect -203 -1045 -191 -1011
rect -283 -1051 -191 -1045
rect -125 -1011 -33 -1005
rect -125 -1045 -113 -1011
rect -45 -1045 -33 -1011
rect -125 -1051 -33 -1045
rect 33 -1011 125 -1005
rect 33 -1045 45 -1011
rect 113 -1045 125 -1011
rect 33 -1051 125 -1045
rect 191 -1011 283 -1005
rect 191 -1045 203 -1011
rect 271 -1045 283 -1011
rect 191 -1051 283 -1045
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 10 l 0.50 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
