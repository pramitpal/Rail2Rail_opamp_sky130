magic
tech sky130A
magscale 1 2
timestamp 1686987678
<< error_p >>
rect -324 -639 -108 -404
rect 108 -639 324 -404
<< mvpdiff >>
rect -258 -527 -174 -470
rect -258 -561 -246 -527
rect -186 -561 -174 -527
rect -258 -573 -174 -561
rect 174 -527 258 -470
rect 174 -561 186 -527
rect 246 -561 258 -527
rect 174 -573 258 -561
<< mvpdiffc >>
rect -246 -561 -186 -527
rect 186 -561 246 -527
<< mvpdiffres >>
rect -258 490 -30 574
rect -258 -470 -174 490
rect -114 -342 -30 490
rect 30 490 258 574
rect 30 -342 114 490
rect -114 -426 114 -342
rect 174 -470 258 490
<< locali >>
rect -262 -561 -246 -527
rect -186 -561 -170 -527
rect 170 -561 186 -527
rect 246 -561 262 -527
<< properties >>
string gencell sky130_fd_pr__res_generic_pd__hv
string library sky130
string parameters w 0.42 l 5 m 1 nx 4 wmin 0.42 lmin 2.10 rho 197 val 11.327k dummy 0 dw 0.02 term 0.0 sterm 0.0 caplen 0.60 snake 1 guard 0 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
