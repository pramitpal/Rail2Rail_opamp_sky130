magic
tech sky130A
timestamp 1681045192
<< error_p >>
rect -87 131 87 133
rect -87 -131 -72 131
rect -54 98 54 100
rect -54 -98 -39 98
rect 39 -98 54 98
rect -54 -100 54 -98
rect 72 -131 87 131
rect -87 -133 87 -131
<< nwell >>
rect -72 -131 72 131
<< mvpmos >>
rect -25 -100 25 100
<< mvpdiff >>
rect -54 94 -25 100
rect -54 -94 -48 94
rect -31 -94 -25 94
rect -54 -100 -25 -94
rect 25 94 54 100
rect 25 -94 31 94
rect 48 -94 54 94
rect 25 -100 54 -94
<< mvpdiffc >>
rect -48 -94 -31 94
rect 31 -94 48 94
<< poly >>
rect -25 100 25 113
rect -25 -113 25 -100
<< locali >>
rect -48 94 -31 102
rect -48 -102 -31 -94
rect 31 94 48 102
rect 31 -102 48 -94
<< viali >>
rect -48 -94 -31 94
rect 31 -94 48 94
<< metal1 >>
rect -51 94 -28 100
rect -51 -94 -48 94
rect -31 -94 -28 94
rect -51 -100 -28 -94
rect 28 94 51 100
rect 28 -94 31 94
rect 48 -94 51 94
rect 28 -100 51 -94
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 2 l 0.50 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
